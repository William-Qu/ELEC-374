library verilog;
use verilog.vl_types.all;
entity TestbenchMultiplier is
end TestbenchMultiplier;
