module RAM (
input clr, clk, write,
input [31:0] dataIn,
input [8:0] Addr,
output [31:0] dataOut
);

reg [31:0] dataOutTemp;

//Make the output value wires
//---------------------------------------------------------------------------------------------------------------------------
wire [31:0]
Mreg0Out, Mreg10Out, Mreg20Out, Mreg30Out, Mreg40Out, Mreg50Out, Mreg60Out, Mreg70Out, Mreg80Out, Mreg90Out,
Mreg1Out, Mreg11Out, Mreg21Out, Mreg31Out, Mreg41Out, Mreg51Out, Mreg61Out, Mreg71Out, Mreg81Out, Mreg91Out,
Mreg2Out, Mreg12Out, Mreg22Out, Mreg32Out, Mreg42Out, Mreg52Out, Mreg62Out, Mreg72Out, Mreg82Out, Mreg92Out,
Mreg3Out, Mreg13Out, Mreg23Out, Mreg33Out, Mreg43Out, Mreg53Out, Mreg63Out, Mreg73Out, Mreg83Out, Mreg93Out,
Mreg4Out, Mreg14Out, Mreg24Out, Mreg34Out, Mreg44Out, Mreg54Out, Mreg64Out, Mreg74Out, Mreg84Out, Mreg94Out,
Mreg5Out, Mreg15Out, Mreg25Out, Mreg35Out, Mreg45Out, Mreg55Out, Mreg65Out, Mreg75Out, Mreg85Out, Mreg95Out,
Mreg6Out, Mreg16Out, Mreg26Out, Mreg36Out, Mreg46Out, Mreg56Out, Mreg66Out, Mreg76Out, Mreg86Out, Mreg96Out, 
Mreg7Out, Mreg17Out, Mreg27Out, Mreg37Out, Mreg47Out, Mreg57Out, Mreg67Out, Mreg77Out, Mreg87Out, Mreg97Out,
Mreg8Out, Mreg18Out, Mreg28Out, Mreg38Out, Mreg48Out, Mreg58Out, Mreg68Out, Mreg78Out, Mreg88Out, Mreg98Out,
Mreg9Out, Mreg19Out, Mreg29Out, Mreg39Out, Mreg49Out, Mreg59Out, Mreg69Out, Mreg79Out, Mreg89Out, Mreg99Out, 
//Hundred Brick
Mreg100Out, Mreg110Out, Mreg120Out, Mreg130Out, Mreg140Out, Mreg150Out, Mreg160Out, Mreg170Out, Mreg180Out, Mreg190Out,
Mreg101Out, Mreg111Out, Mreg121Out, Mreg131Out, Mreg141Out, Mreg151Out, Mreg161Out, Mreg171Out, Mreg181Out, Mreg191Out,
Mreg102Out, Mreg112Out, Mreg122Out, Mreg132Out, Mreg142Out, Mreg152Out, Mreg162Out, Mreg172Out, Mreg182Out, Mreg192Out,
Mreg103Out, Mreg113Out, Mreg123Out, Mreg133Out, Mreg143Out, Mreg153Out, Mreg163Out, Mreg173Out, Mreg183Out, Mreg193Out,
Mreg104Out, Mreg114Out, Mreg124Out, Mreg134Out, Mreg144Out, Mreg154Out, Mreg164Out, Mreg174Out, Mreg184Out, Mreg194Out,
Mreg105Out, Mreg115Out, Mreg125Out, Mreg135Out, Mreg145Out, Mreg155Out, Mreg165Out, Mreg175Out, Mreg185Out, Mreg195Out,
Mreg106Out, Mreg116Out, Mreg126Out, Mreg136Out, Mreg146Out, Mreg156Out, Mreg166Out, Mreg176Out, Mreg186Out, Mreg196Out, 
Mreg107Out, Mreg117Out, Mreg127Out, Mreg137Out, Mreg147Out, Mreg157Out, Mreg167Out, Mreg177Out, Mreg187Out, Mreg197Out,
Mreg108Out, Mreg118Out, Mreg128Out, Mreg138Out, Mreg148Out, Mreg158Out, Mreg168Out, Mreg178Out, Mreg188Out, Mreg198Out,
Mreg109Out, Mreg119Out, Mreg129Out, Mreg139Out, Mreg149Out, Mreg159Out, Mreg169Out, Mreg179Out, Mreg189Out, Mreg199Out, 
//Hundred Brick
Mreg200Out, Mreg210Out, Mreg220Out, Mreg230Out, Mreg240Out, Mreg250Out, Mreg260Out, Mreg270Out, Mreg280Out, Mreg290Out,
Mreg201Out, Mreg211Out, Mreg221Out, Mreg231Out, Mreg241Out, Mreg251Out, Mreg261Out, Mreg271Out, Mreg281Out, Mreg291Out,
Mreg202Out, Mreg212Out, Mreg222Out, Mreg232Out, Mreg242Out, Mreg252Out, Mreg262Out, Mreg272Out, Mreg282Out, Mreg292Out,
Mreg203Out, Mreg213Out, Mreg223Out, Mreg233Out, Mreg243Out, Mreg253Out, Mreg263Out, Mreg273Out, Mreg283Out, Mreg293Out,
Mreg204Out, Mreg214Out, Mreg224Out, Mreg234Out, Mreg244Out, Mreg254Out, Mreg264Out, Mreg274Out, Mreg284Out, Mreg294Out,
Mreg205Out, Mreg215Out, Mreg225Out, Mreg235Out, Mreg245Out, Mreg255Out, Mreg265Out, Mreg275Out, Mreg285Out, Mreg295Out,
Mreg206Out, Mreg216Out, Mreg226Out, Mreg236Out, Mreg246Out, Mreg256Out, Mreg266Out, Mreg276Out, Mreg286Out, Mreg296Out, 
Mreg207Out, Mreg217Out, Mreg227Out, Mreg237Out, Mreg247Out, Mreg257Out, Mreg267Out, Mreg277Out, Mreg287Out, Mreg297Out,
Mreg208Out, Mreg218Out, Mreg228Out, Mreg238Out, Mreg248Out, Mreg258Out, Mreg268Out, Mreg278Out, Mreg288Out, Mreg298Out,
Mreg209Out, Mreg219Out, Mreg229Out, Mreg239Out, Mreg249Out, Mreg259Out, Mreg269Out, Mreg279Out, Mreg289Out, Mreg299Out, 
//Hundred Brick
Mreg300Out, Mreg310Out, Mreg320Out, Mreg330Out, Mreg340Out, Mreg350Out, Mreg360Out, Mreg370Out, Mreg380Out, Mreg390Out,
Mreg301Out, Mreg311Out, Mreg321Out, Mreg331Out, Mreg341Out, Mreg351Out, Mreg361Out, Mreg371Out, Mreg381Out, Mreg391Out,
Mreg302Out, Mreg312Out, Mreg322Out, Mreg332Out, Mreg342Out, Mreg352Out, Mreg362Out, Mreg372Out, Mreg382Out, Mreg392Out,
Mreg303Out, Mreg313Out, Mreg323Out, Mreg333Out, Mreg343Out, Mreg353Out, Mreg363Out, Mreg373Out, Mreg383Out, Mreg393Out,
Mreg304Out, Mreg314Out, Mreg324Out, Mreg334Out, Mreg344Out, Mreg354Out, Mreg364Out, Mreg374Out, Mreg384Out, Mreg394Out,
Mreg305Out, Mreg315Out, Mreg325Out, Mreg335Out, Mreg345Out, Mreg355Out, Mreg365Out, Mreg375Out, Mreg385Out, Mreg395Out,
Mreg306Out, Mreg316Out, Mreg326Out, Mreg336Out, Mreg346Out, Mreg356Out, Mreg366Out, Mreg376Out, Mreg386Out, Mreg396Out, 
Mreg307Out, Mreg317Out, Mreg327Out, Mreg337Out, Mreg347Out, Mreg357Out, Mreg367Out, Mreg377Out, Mreg387Out, Mreg397Out,
Mreg308Out, Mreg318Out, Mreg328Out, Mreg338Out, Mreg348Out, Mreg358Out, Mreg368Out, Mreg378Out, Mreg388Out, Mreg398Out,
Mreg309Out, Mreg319Out, Mreg329Out, Mreg339Out, Mreg349Out, Mreg359Out, Mreg369Out, Mreg379Out, Mreg389Out, Mreg399Out, 
//Hundred Brick
Mreg400Out, Mreg410Out, Mreg420Out, Mreg430Out, Mreg440Out, Mreg450Out, Mreg460Out, Mreg470Out, Mreg480Out, Mreg490Out,
Mreg401Out, Mreg411Out, Mreg421Out, Mreg431Out, Mreg441Out, Mreg451Out, Mreg461Out, Mreg471Out, Mreg481Out, Mreg491Out,
Mreg402Out, Mreg412Out, Mreg422Out, Mreg432Out, Mreg442Out, Mreg452Out, Mreg462Out, Mreg472Out, Mreg482Out, Mreg492Out,
Mreg403Out, Mreg413Out, Mreg423Out, Mreg433Out, Mreg443Out, Mreg453Out, Mreg463Out, Mreg473Out, Mreg483Out, Mreg493Out,
Mreg404Out, Mreg414Out, Mreg424Out, Mreg434Out, Mreg444Out, Mreg454Out, Mreg464Out, Mreg474Out, Mreg484Out, Mreg494Out,
Mreg405Out, Mreg415Out, Mreg425Out, Mreg435Out, Mreg445Out, Mreg455Out, Mreg465Out, Mreg475Out, Mreg485Out, Mreg495Out,
Mreg406Out, Mreg416Out, Mreg426Out, Mreg436Out, Mreg446Out, Mreg456Out, Mreg466Out, Mreg476Out, Mreg486Out, Mreg496Out, 
Mreg407Out, Mreg417Out, Mreg427Out, Mreg437Out, Mreg447Out, Mreg457Out, Mreg467Out, Mreg477Out, Mreg487Out, Mreg497Out,
Mreg408Out, Mreg418Out, Mreg428Out, Mreg438Out, Mreg448Out, Mreg458Out, Mreg468Out, Mreg478Out, Mreg488Out, Mreg498Out,
Mreg409Out, Mreg419Out, Mreg429Out, Mreg439Out, Mreg449Out, Mreg459Out, Mreg469Out, Mreg479Out, Mreg489Out, Mreg499Out, 
//Hundred Brick
Mreg500Out, Mreg501Out, Mreg502Out, Mreg503Out, Mreg504Out, Mreg505Out, Mreg506Out, Mreg507Out, Mreg508Out, Mreg509Out, 
Mreg510Out, Mreg511Out;
//---------------------------------------------------------------------------------------------------------------------------
//Finish making the output value wires

//Make the input enable signals 
//---------------------------------------------------------------------------------------------------------------------------
reg [31:0]
Mreg0Ins, Mreg10Ins, Mreg20Ins, Mreg30Ins, Mreg40Ins, Mreg50Ins, Mreg60Ins, Mreg70Ins, Mreg80Ins, Mreg90Ins,
Mreg1Ins, Mreg11Ins, Mreg21Ins, Mreg31Ins, Mreg41Ins, Mreg51Ins, Mreg61Ins, Mreg71Ins, Mreg81Ins, Mreg91Ins,
Mreg2Ins, Mreg12Ins, Mreg22Ins, Mreg32Ins, Mreg42Ins, Mreg52Ins, Mreg62Ins, Mreg72Ins, Mreg82Ins, Mreg92Ins,
Mreg3Ins, Mreg13Ins, Mreg23Ins, Mreg33Ins, Mreg43Ins, Mreg53Ins, Mreg63Ins, Mreg73Ins, Mreg83Ins, Mreg93Ins,
Mreg4Ins, Mreg14Ins, Mreg24Ins, Mreg34Ins, Mreg44Ins, Mreg54Ins, Mreg64Ins, Mreg74Ins, Mreg84Ins, Mreg94Ins,
Mreg5Ins, Mreg15Ins, Mreg25Ins, Mreg35Ins, Mreg45Ins, Mreg55Ins, Mreg65Ins, Mreg75Ins, Mreg85Ins, Mreg95Ins,
Mreg6Ins, Mreg16Ins, Mreg26Ins, Mreg36Ins, Mreg46Ins, Mreg56Ins, Mreg66Ins, Mreg76Ins, Mreg86Ins, Mreg96Ins, 
Mreg7Ins, Mreg17Ins, Mreg27Ins, Mreg37Ins, Mreg47Ins, Mreg57Ins, Mreg67Ins, Mreg77Ins, Mreg87Ins, Mreg97Ins,
Mreg8Ins, Mreg18Ins, Mreg28Ins, Mreg38Ins, Mreg48Ins, Mreg58Ins, Mreg68Ins, Mreg78Ins, Mreg88Ins, Mreg98Ins,
Mreg9Ins, Mreg19Ins, Mreg29Ins, Mreg39Ins, Mreg49Ins, Mreg59Ins, Mreg69Ins, Mreg79Ins, Mreg89Ins, Mreg99Ins, 
//Hundred Brick
Mreg100Ins, Mreg110Ins, Mreg120Ins, Mreg130Ins, Mreg140Ins, Mreg150Ins, Mreg160Ins, Mreg170Ins, Mreg180Ins, Mreg190Ins,
Mreg101Ins, Mreg111Ins, Mreg121Ins, Mreg131Ins, Mreg141Ins, Mreg151Ins, Mreg161Ins, Mreg171Ins, Mreg181Ins, Mreg191Ins,
Mreg102Ins, Mreg112Ins, Mreg122Ins, Mreg132Ins, Mreg142Ins, Mreg152Ins, Mreg162Ins, Mreg172Ins, Mreg182Ins, Mreg192Ins,
Mreg103Ins, Mreg113Ins, Mreg123Ins, Mreg133Ins, Mreg143Ins, Mreg153Ins, Mreg163Ins, Mreg173Ins, Mreg183Ins, Mreg193Ins,
Mreg104Ins, Mreg114Ins, Mreg124Ins, Mreg134Ins, Mreg144Ins, Mreg154Ins, Mreg164Ins, Mreg174Ins, Mreg184Ins, Mreg194Ins,
Mreg105Ins, Mreg115Ins, Mreg125Ins, Mreg135Ins, Mreg145Ins, Mreg155Ins, Mreg165Ins, Mreg175Ins, Mreg185Ins, Mreg195Ins,
Mreg106Ins, Mreg116Ins, Mreg126Ins, Mreg136Ins, Mreg146Ins, Mreg156Ins, Mreg166Ins, Mreg176Ins, Mreg186Ins, Mreg196Ins, 
Mreg107Ins, Mreg117Ins, Mreg127Ins, Mreg137Ins, Mreg147Ins, Mreg157Ins, Mreg167Ins, Mreg177Ins, Mreg187Ins, Mreg197Ins,
Mreg108Ins, Mreg118Ins, Mreg128Ins, Mreg138Ins, Mreg148Ins, Mreg158Ins, Mreg168Ins, Mreg178Ins, Mreg188Ins, Mreg198Ins,
Mreg109Ins, Mreg119Ins, Mreg129Ins, Mreg139Ins, Mreg149Ins, Mreg159Ins, Mreg169Ins, Mreg179Ins, Mreg189Ins, Mreg199Ins, 
//Hundred Brick 
Mreg200Ins, Mreg210Ins, Mreg220Ins, Mreg230Ins, Mreg240Ins, Mreg250Ins, Mreg260Ins, Mreg270Ins, Mreg280Ins, Mreg290Ins,
Mreg201Ins, Mreg211Ins, Mreg221Ins, Mreg231Ins, Mreg241Ins, Mreg251Ins, Mreg261Ins, Mreg271Ins, Mreg281Ins, Mreg291Ins,
Mreg202Ins, Mreg212Ins, Mreg222Ins, Mreg232Ins, Mreg242Ins, Mreg252Ins, Mreg262Ins, Mreg272Ins, Mreg282Ins, Mreg292Ins,
Mreg203Ins, Mreg213Ins, Mreg223Ins, Mreg233Ins, Mreg243Ins, Mreg253Ins, Mreg263Ins, Mreg273Ins, Mreg283Ins, Mreg293Ins,
Mreg204Ins, Mreg214Ins, Mreg224Ins, Mreg234Ins, Mreg244Ins, Mreg254Ins, Mreg264Ins, Mreg274Ins, Mreg284Ins, Mreg294Ins,
Mreg205Ins, Mreg215Ins, Mreg225Ins, Mreg235Ins, Mreg245Ins, Mreg255Ins, Mreg265Ins, Mreg275Ins, Mreg285Ins, Mreg295Ins,
Mreg206Ins, Mreg216Ins, Mreg226Ins, Mreg236Ins, Mreg246Ins, Mreg256Ins, Mreg266Ins, Mreg276Ins, Mreg286Ins, Mreg296Ins, 
Mreg207Ins, Mreg217Ins, Mreg227Ins, Mreg237Ins, Mreg247Ins, Mreg257Ins, Mreg267Ins, Mreg277Ins, Mreg287Ins, Mreg297Ins,
Mreg208Ins, Mreg218Ins, Mreg228Ins, Mreg238Ins, Mreg248Ins, Mreg258Ins, Mreg268Ins, Mreg278Ins, Mreg288Ins, Mreg298Ins,
Mreg209Ins, Mreg219Ins, Mreg229Ins, Mreg239Ins, Mreg249Ins, Mreg259Ins, Mreg269Ins, Mreg279Ins, Mreg289Ins, Mreg299Ins, 
//Hundred Brick  
Mreg300Ins, Mreg310Ins, Mreg320Ins, Mreg330Ins, Mreg340Ins, Mreg350Ins, Mreg360Ins, Mreg370Ins, Mreg380Ins, Mreg390Ins,
Mreg301Ins, Mreg311Ins, Mreg321Ins, Mreg331Ins, Mreg341Ins, Mreg351Ins, Mreg361Ins, Mreg371Ins, Mreg381Ins, Mreg391Ins,
Mreg302Ins, Mreg312Ins, Mreg322Ins, Mreg332Ins, Mreg342Ins, Mreg352Ins, Mreg362Ins, Mreg372Ins, Mreg382Ins, Mreg392Ins,
Mreg303Ins, Mreg313Ins, Mreg323Ins, Mreg333Ins, Mreg343Ins, Mreg353Ins, Mreg363Ins, Mreg373Ins, Mreg383Ins, Mreg393Ins,
Mreg304Ins, Mreg314Ins, Mreg324Ins, Mreg334Ins, Mreg344Ins, Mreg354Ins, Mreg364Ins, Mreg374Ins, Mreg384Ins, Mreg394Ins,
Mreg305Ins, Mreg315Ins, Mreg325Ins, Mreg335Ins, Mreg345Ins, Mreg355Ins, Mreg365Ins, Mreg375Ins, Mreg385Ins, Mreg395Ins,
Mreg306Ins, Mreg316Ins, Mreg326Ins, Mreg336Ins, Mreg346Ins, Mreg356Ins, Mreg366Ins, Mreg376Ins, Mreg386Ins, Mreg396Ins, 
Mreg307Ins, Mreg317Ins, Mreg327Ins, Mreg337Ins, Mreg347Ins, Mreg357Ins, Mreg367Ins, Mreg377Ins, Mreg387Ins, Mreg397Ins,
Mreg308Ins, Mreg318Ins, Mreg328Ins, Mreg338Ins, Mreg348Ins, Mreg358Ins, Mreg368Ins, Mreg378Ins, Mreg388Ins, Mreg398Ins,
Mreg309Ins, Mreg319Ins, Mreg329Ins, Mreg339Ins, Mreg349Ins, Mreg359Ins, Mreg369Ins, Mreg379Ins, Mreg389Ins, Mreg399Ins, 
//Hundred Brick   
Mreg400Ins, Mreg410Ins, Mreg420Ins, Mreg430Ins, Mreg440Ins, Mreg450Ins, Mreg460Ins, Mreg470Ins, Mreg480Ins, Mreg490Ins,
Mreg401Ins, Mreg411Ins, Mreg421Ins, Mreg431Ins, Mreg441Ins, Mreg451Ins, Mreg461Ins, Mreg471Ins, Mreg481Ins, Mreg491Ins,
Mreg402Ins, Mreg412Ins, Mreg422Ins, Mreg432Ins, Mreg442Ins, Mreg452Ins, Mreg462Ins, Mreg472Ins, Mreg482Ins, Mreg492Ins,
Mreg403Ins, Mreg413Ins, Mreg423Ins, Mreg433Ins, Mreg443Ins, Mreg453Ins, Mreg463Ins, Mreg473Ins, Mreg483Ins, Mreg493Ins,
Mreg404Ins, Mreg414Ins, Mreg424Ins, Mreg434Ins, Mreg444Ins, Mreg454Ins, Mreg464Ins, Mreg474Ins, Mreg484Ins, Mreg494Ins,
Mreg405Ins, Mreg415Ins, Mreg425Ins, Mreg435Ins, Mreg445Ins, Mreg455Ins, Mreg465Ins, Mreg475Ins, Mreg485Ins, Mreg495Ins,
Mreg406Ins, Mreg416Ins, Mreg426Ins, Mreg436Ins, Mreg446Ins, Mreg456Ins, Mreg466Ins, Mreg476Ins, Mreg486Ins, Mreg496Ins, 
Mreg407Ins, Mreg417Ins, Mreg427Ins, Mreg437Ins, Mreg447Ins, Mreg457Ins, Mreg467Ins, Mreg477Ins, Mreg487Ins, Mreg497Ins,
Mreg408Ins, Mreg418Ins, Mreg428Ins, Mreg438Ins, Mreg448Ins, Mreg458Ins, Mreg468Ins, Mreg478Ins, Mreg488Ins, Mreg498Ins,
Mreg409Ins, Mreg419Ins, Mreg429Ins, Mreg439Ins, Mreg449Ins, Mreg459Ins, Mreg469Ins, Mreg479Ins, Mreg489Ins, Mreg499Ins, 
//Hundred Brick  
Mreg500Ins, Mreg501Ins, Mreg502Ins, Mreg503Ins, Mreg504Ins, Mreg505Ins, Mreg506Ins, Mreg507Ins, Mreg508Ins, Mreg509Ins, 
Mreg510Ins, Mreg511Ins;
//---------------------------------------------------------------------------------------------------------------------------
//Finish making the input enable signals

	//Generate the 512 32-bit registers
	generate
		reg32bit Mreg0  (Mreg0Out,  dataIn, clr, clk, Mreg0Ins);
		reg32bit Mreg1  (Mreg1Out,  dataIn, clr, clk, Mreg1Ins);
		reg32bit Mreg2  (Mreg2Out,  dataIn, clr, clk, Mreg2Ins);
		reg32bit Mreg3  (Mreg3Out,  dataIn, clr, clk, Mreg3Ins);
		reg32bit Mreg4  (Mreg4Out,  dataIn, clr, clk, Mreg4Ins);
		reg32bit Mreg5  (Mreg5Out,  dataIn, clr, clk, Mreg5Ins);
		reg32bit Mreg6  (Mreg6Out,  dataIn, clr, clk, Mreg6Ins);
		reg32bit Mreg7  (Mreg7Out,  dataIn, clr, clk, Mreg7Ins);
		reg32bit Mreg8  (Mreg8Out,  dataIn, clr, clk, Mreg8Ins);
		reg32bit Mreg9  (Mreg9Out,  dataIn, clr, clk, Mreg9Ins);
		reg32bit Mreg10 (Mreg10Out, dataIn, clr, clk, Mreg10Ins);
		reg32bit Mreg11 (Mreg11Out, dataIn, clr, clk, Mreg11Ins);
		reg32bit Mreg12 (Mreg12Out, dataIn, clr, clk, Mreg12Ins);
		reg32bit Mreg13 (Mreg13Out, dataIn, clr, clk, Mreg13Ins);
		reg32bit Mreg14 (Mreg14Out, dataIn, clr, clk, Mreg14Ins);
		reg32bit Mreg15 (Mreg15Out, dataIn, clr, clk, Mreg15Ins);
		reg32bit Mreg16 (Mreg16Out, dataIn, clr, clk, Mreg16Ins);
		reg32bit Mreg17 (Mreg17Out, dataIn, clr, clk, Mreg17Ins);
		reg32bit Mreg18 (Mreg18Out, dataIn, clr, clk, Mreg18Ins);
		reg32bit Mreg19 (Mreg19Out, dataIn, clr, clk, Mreg19Ins);
		reg32bit Mreg20 (Mreg20Out, dataIn, clr, clk, Mreg20Ins);
		reg32bit Mreg21 (Mreg21Out, dataIn, clr, clk, Mreg21Ins);
		reg32bit Mreg22 (Mreg22Out, dataIn, clr, clk, Mreg22Ins);
		reg32bit Mreg23 (Mreg23Out, dataIn, clr, clk, Mreg23Ins);
		reg32bit Mreg24 (Mreg24Out, dataIn, clr, clk, Mreg24Ins);
		reg32bit Mreg25 (Mreg25Out, dataIn, clr, clk, Mreg25Ins);
		reg32bit Mreg26 (Mreg26Out, dataIn, clr, clk, Mreg26Ins);
		reg32bit Mreg27 (Mreg27Out, dataIn, clr, clk, Mreg27Ins);
		reg32bit Mreg28 (Mreg28Out, dataIn, clr, clk, Mreg28Ins);
		reg32bit Mreg29 (Mreg29Out, dataIn, clr, clk, Mreg29Ins);
		reg32bit Mreg30 (Mreg30Out, dataIn, clr, clk, Mreg30Ins);
		reg32bit Mreg31 (Mreg31Out, dataIn, clr, clk, Mreg31Ins);
		reg32bit Mreg32 (Mreg32Out, dataIn, clr, clk, Mreg32Ins);
		reg32bit Mreg33 (Mreg33Out, dataIn, clr, clk, Mreg33Ins);
		reg32bit Mreg34 (Mreg34Out, dataIn, clr, clk, Mreg34Ins);
		reg32bit Mreg35 (Mreg35Out, dataIn, clr, clk, Mreg35Ins);
		reg32bit Mreg36 (Mreg36Out, dataIn, clr, clk, Mreg36Ins);
		reg32bit Mreg37 (Mreg37Out, dataIn, clr, clk, Mreg37Ins);
		reg32bit Mreg38 (Mreg38Out, dataIn, clr, clk, Mreg38Ins);
		reg32bit Mreg39 (Mreg39Out, dataIn, clr, clk, Mreg39Ins);
		reg32bit Mreg40 (Mreg40Out, dataIn, clr, clk, Mreg40Ins);
		reg32bit Mreg41 (Mreg41Out, dataIn, clr, clk, Mreg41Ins);
		reg32bit Mreg42 (Mreg42Out, dataIn, clr, clk, Mreg42Ins);
		reg32bit Mreg43 (Mreg43Out, dataIn, clr, clk, Mreg43Ins);
		reg32bit Mreg44 (Mreg44Out, dataIn, clr, clk, Mreg44Ins);
		reg32bit Mreg45 (Mreg45Out, dataIn, clr, clk, Mreg45Ins);
		reg32bit Mreg46 (Mreg46Out, dataIn, clr, clk, Mreg46Ins);
		reg32bit Mreg47 (Mreg47Out, dataIn, clr, clk, Mreg47Ins);
		reg32bit Mreg48 (Mreg48Out, dataIn, clr, clk, Mreg48Ins);
		reg32bit Mreg49 (Mreg49Out, dataIn, clr, clk, Mreg49Ins);
		reg32bit Mreg50 (Mreg50Out, dataIn, clr, clk, Mreg50Ins);
		reg32bit Mreg51 (Mreg51Out, dataIn, clr, clk, Mreg51Ins);
		reg32bit Mreg52 (Mreg52Out, dataIn, clr, clk, Mreg52Ins);
		reg32bit Mreg53 (Mreg53Out, dataIn, clr, clk, Mreg53Ins);
		reg32bit Mreg54 (Mreg54Out, dataIn, clr, clk, Mreg54Ins);
		reg32bit Mreg55 (Mreg55Out, dataIn, clr, clk, Mreg55Ins);
		reg32bit Mreg56 (Mreg56Out, dataIn, clr, clk, Mreg56Ins);
		reg32bit Mreg57 (Mreg57Out, dataIn, clr, clk, Mreg57Ins);
		reg32bit Mreg58 (Mreg58Out, dataIn, clr, clk, Mreg58Ins);
		reg32bit Mreg59 (Mreg59Out, dataIn, clr, clk, Mreg59Ins);
		reg32bit Mreg60 (Mreg60Out, dataIn, clr, clk, Mreg60Ins);
		reg32bit Mreg61 (Mreg61Out, dataIn, clr, clk, Mreg61Ins);
		reg32bit Mreg62 (Mreg62Out, dataIn, clr, clk, Mreg62Ins);
		reg32bit Mreg63 (Mreg63Out, dataIn, clr, clk, Mreg63Ins);
		reg32bit Mreg64 (Mreg64Out, dataIn, clr, clk, Mreg64Ins);
		reg32bit Mreg65 (Mreg65Out, dataIn, clr, clk, Mreg65Ins);
		reg32bit Mreg66 (Mreg66Out, dataIn, clr, clk, Mreg66Ins);
		reg32bit Mreg67 (Mreg67Out, dataIn, clr, clk, Mreg67Ins);
		reg32bit Mreg68 (Mreg68Out, dataIn, clr, clk, Mreg68Ins);
		reg32bit Mreg69 (Mreg69Out, dataIn, clr, clk, Mreg69Ins);
		reg32bit Mreg70 (Mreg70Out, dataIn, clr, clk, Mreg70Ins);
		reg32bit Mreg71 (Mreg71Out, dataIn, clr, clk, Mreg71Ins);
		reg32bit Mreg72 (Mreg72Out, dataIn, clr, clk, Mreg72Ins);
		reg32bit Mreg73 (Mreg73Out, dataIn, clr, clk, Mreg73Ins);
		reg32bit Mreg74 (Mreg74Out, dataIn, clr, clk, Mreg74Ins);
		reg32bit Mreg75 (Mreg75Out, dataIn, clr, clk, Mreg75Ins);
		reg32bit Mreg76 (Mreg76Out, dataIn, clr, clk, Mreg76Ins);
		reg32bit Mreg77 (Mreg77Out, dataIn, clr, clk, Mreg77Ins);
		reg32bit Mreg78 (Mreg78Out, dataIn, clr, clk, Mreg78Ins);
		reg32bit Mreg79 (Mreg79Out, dataIn, clr, clk, Mreg79Ins);
		reg32bit Mreg80 (Mreg80Out, dataIn, clr, clk, Mreg80Ins);
		reg32bit Mreg81 (Mreg81Out, dataIn, clr, clk, Mreg81Ins);
		reg32bit Mreg82 (Mreg82Out, dataIn, clr, clk, Mreg82Ins);
		reg32bit Mreg83 (Mreg83Out, dataIn, clr, clk, Mreg83Ins);
		reg32bit Mreg84 (Mreg84Out, dataIn, clr, clk, Mreg84Ins);
		reg32bit Mreg85 (Mreg85Out, dataIn, clr, clk, Mreg85Ins);
		reg32bit Mreg86 (Mreg86Out, dataIn, clr, clk, Mreg86Ins);
		reg32bit Mreg87 (Mreg87Out, dataIn, clr, clk, Mreg87Ins);
		reg32bit Mreg88 (Mreg88Out, dataIn, clr, clk, Mreg88Ins);
		reg32bit Mreg89 (Mreg89Out, dataIn, clr, clk, Mreg89Ins);
		reg32bit Mreg90 (Mreg90Out, dataIn, clr, clk, Mreg90Ins);
		reg32bit Mreg91 (Mreg91Out, dataIn, clr, clk, Mreg91Ins);
		reg32bit Mreg92 (Mreg92Out, dataIn, clr, clk, Mreg92Ins);
		reg32bit Mreg93 (Mreg93Out, dataIn, clr, clk, Mreg93Ins);
		reg32bit Mreg94 (Mreg94Out, dataIn, clr, clk, Mreg94Ins);
		reg32bit Mreg95 (Mreg95Out, dataIn, clr, clk, Mreg95Ins);
		reg32bit Mreg96 (Mreg96Out, dataIn, clr, clk, Mreg96Ins);
		reg32bit Mreg97 (Mreg97Out, dataIn, clr, clk, Mreg97Ins);
		reg32bit Mreg98 (Mreg98Out, dataIn, clr, clk, Mreg98Ins);
		reg32bit Mreg99 (Mreg99Out, dataIn, clr, clk, Mreg99Ins);
		//Break for a hundred
		reg32bit Mreg100 (Mreg100Out, dataIn, clr, clk, Mreg100Ins);
		reg32bit Mreg101 (Mreg101Out, dataIn, clr, clk, Mreg101Ins);
		reg32bit Mreg102 (Mreg102Out, dataIn, clr, clk, Mreg102Ins);
		reg32bit Mreg103 (Mreg103Out, dataIn, clr, clk, Mreg103Ins);
		reg32bit Mreg104 (Mreg104Out, dataIn, clr, clk, Mreg104Ins);
		reg32bit Mreg105 (Mreg105Out, dataIn, clr, clk, Mreg105Ins);
		reg32bit Mreg106 (Mreg106Out, dataIn, clr, clk, Mreg106Ins);
		reg32bit Mreg107 (Mreg107Out, dataIn, clr, clk, Mreg107Ins);
		reg32bit Mreg108 (Mreg108Out, dataIn, clr, clk, Mreg108Ins);
		reg32bit Mreg109 (Mreg109Out, dataIn, clr, clk, Mreg109Ins);
		reg32bit Mreg110 (Mreg110Out, dataIn, clr, clk, Mreg110Ins);
		reg32bit Mreg111 (Mreg111Out, dataIn, clr, clk, Mreg111Ins);
		reg32bit Mreg112 (Mreg112Out, dataIn, clr, clk, Mreg112Ins);
		reg32bit Mreg113 (Mreg113Out, dataIn, clr, clk, Mreg113Ins);
		reg32bit Mreg114 (Mreg114Out, dataIn, clr, clk, Mreg114Ins);
		reg32bit Mreg115 (Mreg115Out, dataIn, clr, clk, Mreg115Ins);
		reg32bit Mreg116 (Mreg116Out, dataIn, clr, clk, Mreg116Ins);
		reg32bit Mreg117 (Mreg117Out, dataIn, clr, clk, Mreg117Ins);
		reg32bit Mreg118 (Mreg118Out, dataIn, clr, clk, Mreg118Ins);
		reg32bit Mreg119 (Mreg119Out, dataIn, clr, clk, Mreg119Ins);
		reg32bit Mreg120 (Mreg120Out, dataIn, clr, clk, Mreg120Ins);
		reg32bit Mreg121 (Mreg121Out, dataIn, clr, clk, Mreg121Ins);
		reg32bit Mreg122 (Mreg122Out, dataIn, clr, clk, Mreg122Ins);
		reg32bit Mreg123 (Mreg123Out, dataIn, clr, clk, Mreg123Ins);
		reg32bit Mreg124 (Mreg124Out, dataIn, clr, clk, Mreg124Ins);
		reg32bit Mreg125 (Mreg125Out, dataIn, clr, clk, Mreg125Ins);
		reg32bit Mreg126 (Mreg126Out, dataIn, clr, clk, Mreg126Ins);
		reg32bit Mreg127 (Mreg127Out, dataIn, clr, clk, Mreg127Ins);
		reg32bit Mreg128 (Mreg128Out, dataIn, clr, clk, Mreg128Ins);
		reg32bit Mreg129 (Mreg129Out, dataIn, clr, clk, Mreg129Ins);
		reg32bit Mreg130 (Mreg130Out, dataIn, clr, clk, Mreg130Ins);
		reg32bit Mreg131 (Mreg131Out, dataIn, clr, clk, Mreg131Ins);
		reg32bit Mreg132 (Mreg132Out, dataIn, clr, clk, Mreg132Ins);
		reg32bit Mreg133 (Mreg133Out, dataIn, clr, clk, Mreg133Ins);
		reg32bit Mreg134 (Mreg134Out, dataIn, clr, clk, Mreg134Ins);
		reg32bit Mreg135 (Mreg135Out, dataIn, clr, clk, Mreg135Ins);
		reg32bit Mreg136 (Mreg136Out, dataIn, clr, clk, Mreg136Ins);
		reg32bit Mreg137 (Mreg137Out, dataIn, clr, clk, Mreg137Ins);
		reg32bit Mreg138 (Mreg138Out, dataIn, clr, clk, Mreg138Ins);
		reg32bit Mreg139 (Mreg139Out, dataIn, clr, clk, Mreg139Ins);
		reg32bit Mreg140 (Mreg140Out, dataIn, clr, clk, Mreg140Ins);
		reg32bit Mreg141 (Mreg141Out, dataIn, clr, clk, Mreg141Ins);
		reg32bit Mreg142 (Mreg142Out, dataIn, clr, clk, Mreg142Ins);
		reg32bit Mreg143 (Mreg143Out, dataIn, clr, clk, Mreg143Ins);
		reg32bit Mreg144 (Mreg144Out, dataIn, clr, clk, Mreg144Ins);
		reg32bit Mreg145 (Mreg145Out, dataIn, clr, clk, Mreg145Ins);
		reg32bit Mreg146 (Mreg146Out, dataIn, clr, clk, Mreg146Ins);
		reg32bit Mreg147 (Mreg147Out, dataIn, clr, clk, Mreg147Ins);
		reg32bit Mreg148 (Mreg148Out, dataIn, clr, clk, Mreg148Ins);
		reg32bit Mreg149 (Mreg149Out, dataIn, clr, clk, Mreg149Ins);
		reg32bit Mreg150 (Mreg150Out, dataIn, clr, clk, Mreg150Ins);
		reg32bit Mreg151 (Mreg151Out, dataIn, clr, clk, Mreg151Ins);
		reg32bit Mreg152 (Mreg152Out, dataIn, clr, clk, Mreg152Ins);
		reg32bit Mreg153 (Mreg153Out, dataIn, clr, clk, Mreg153Ins);
		reg32bit Mreg154 (Mreg154Out, dataIn, clr, clk, Mreg154Ins);
		reg32bit Mreg155 (Mreg155Out, dataIn, clr, clk, Mreg155Ins);
		reg32bit Mreg156 (Mreg156Out, dataIn, clr, clk, Mreg156Ins);
		reg32bit Mreg157 (Mreg157Out, dataIn, clr, clk, Mreg157Ins);
		reg32bit Mreg158 (Mreg158Out, dataIn, clr, clk, Mreg158Ins);
		reg32bit Mreg159 (Mreg159Out, dataIn, clr, clk, Mreg159Ins);
		reg32bit Mreg160 (Mreg160Out, dataIn, clr, clk, Mreg160Ins);
		reg32bit Mreg161 (Mreg161Out, dataIn, clr, clk, Mreg161Ins);
		reg32bit Mreg162 (Mreg162Out, dataIn, clr, clk, Mreg162Ins);
		reg32bit Mreg163 (Mreg163Out, dataIn, clr, clk, Mreg163Ins);
		reg32bit Mreg164 (Mreg164Out, dataIn, clr, clk, Mreg164Ins);
		reg32bit Mreg165 (Mreg165Out, dataIn, clr, clk, Mreg165Ins);
		reg32bit Mreg166 (Mreg166Out, dataIn, clr, clk, Mreg166Ins);
		reg32bit Mreg167 (Mreg167Out, dataIn, clr, clk, Mreg167Ins);
		reg32bit Mreg168 (Mreg168Out, dataIn, clr, clk, Mreg168Ins);
		reg32bit Mreg169 (Mreg169Out, dataIn, clr, clk, Mreg169Ins);
		reg32bit Mreg170 (Mreg170Out, dataIn, clr, clk, Mreg170Ins);
		reg32bit Mreg171 (Mreg171Out, dataIn, clr, clk, Mreg171Ins);
		reg32bit Mreg172 (Mreg172Out, dataIn, clr, clk, Mreg172Ins);
		reg32bit Mreg173 (Mreg173Out, dataIn, clr, clk, Mreg173Ins);
		reg32bit Mreg174 (Mreg174Out, dataIn, clr, clk, Mreg174Ins);
		reg32bit Mreg175 (Mreg175Out, dataIn, clr, clk, Mreg175Ins);
		reg32bit Mreg176 (Mreg176Out, dataIn, clr, clk, Mreg176Ins);
		reg32bit Mreg177 (Mreg177Out, dataIn, clr, clk, Mreg177Ins);
		reg32bit Mreg178 (Mreg178Out, dataIn, clr, clk, Mreg178Ins);
		reg32bit Mreg179 (Mreg179Out, dataIn, clr, clk, Mreg179Ins);
		reg32bit Mreg180 (Mreg180Out, dataIn, clr, clk, Mreg180Ins);
		reg32bit Mreg181 (Mreg181Out, dataIn, clr, clk, Mreg181Ins);
		reg32bit Mreg182 (Mreg182Out, dataIn, clr, clk, Mreg182Ins);
		reg32bit Mreg183 (Mreg183Out, dataIn, clr, clk, Mreg183Ins);
		reg32bit Mreg184 (Mreg184Out, dataIn, clr, clk, Mreg184Ins);
		reg32bit Mreg185 (Mreg185Out, dataIn, clr, clk, Mreg185Ins);
		reg32bit Mreg186 (Mreg186Out, dataIn, clr, clk, Mreg186Ins);
		reg32bit Mreg187 (Mreg187Out, dataIn, clr, clk, Mreg187Ins);
		reg32bit Mreg188 (Mreg188Out, dataIn, clr, clk, Mreg188Ins);
		reg32bit Mreg189 (Mreg189Out, dataIn, clr, clk, Mreg189Ins);
		reg32bit Mreg190 (Mreg190Out, dataIn, clr, clk, Mreg190Ins);
		reg32bit Mreg191 (Mreg191Out, dataIn, clr, clk, Mreg191Ins);
		reg32bit Mreg192 (Mreg192Out, dataIn, clr, clk, Mreg192Ins);
		reg32bit Mreg193 (Mreg193Out, dataIn, clr, clk, Mreg193Ins);
		reg32bit Mreg194 (Mreg194Out, dataIn, clr, clk, Mreg194Ins);
		reg32bit Mreg195 (Mreg195Out, dataIn, clr, clk, Mreg195Ins);
		reg32bit Mreg196 (Mreg196Out, dataIn, clr, clk, Mreg196Ins);
		reg32bit Mreg197 (Mreg197Out, dataIn, clr, clk, Mreg197Ins);
		reg32bit Mreg198 (Mreg198Out, dataIn, clr, clk, Mreg198Ins);
		reg32bit Mreg199 (Mreg199Out, dataIn, clr, clk, Mreg199Ins);
		//Break for a hundred
		reg32bit Mreg200 (Mreg200Out, dataIn, clr, clk, Mreg200Ins);
		reg32bit Mreg201 (Mreg201Out, dataIn, clr, clk, Mreg201Ins);
		reg32bit Mreg202 (Mreg202Out, dataIn, clr, clk, Mreg202Ins);
		reg32bit Mreg203 (Mreg203Out, dataIn, clr, clk, Mreg203Ins);
		reg32bit Mreg204 (Mreg204Out, dataIn, clr, clk, Mreg204Ins);
		reg32bit Mreg205 (Mreg205Out, dataIn, clr, clk, Mreg205Ins);
		reg32bit Mreg206 (Mreg206Out, dataIn, clr, clk, Mreg206Ins);
		reg32bit Mreg207 (Mreg207Out, dataIn, clr, clk, Mreg207Ins);
		reg32bit Mreg208 (Mreg208Out, dataIn, clr, clk, Mreg208Ins);
		reg32bit Mreg209 (Mreg209Out, dataIn, clr, clk, Mreg209Ins);
		reg32bit Mreg210 (Mreg210Out, dataIn, clr, clk, Mreg210Ins);
		reg32bit Mreg211 (Mreg211Out, dataIn, clr, clk, Mreg211Ins);
		reg32bit Mreg212 (Mreg212Out, dataIn, clr, clk, Mreg212Ins);
		reg32bit Mreg213 (Mreg213Out, dataIn, clr, clk, Mreg213Ins);
		reg32bit Mreg214 (Mreg214Out, dataIn, clr, clk, Mreg214Ins);
		reg32bit Mreg215 (Mreg215Out, dataIn, clr, clk, Mreg215Ins);
		reg32bit Mreg216 (Mreg216Out, dataIn, clr, clk, Mreg216Ins);
		reg32bit Mreg217 (Mreg217Out, dataIn, clr, clk, Mreg217Ins);
		reg32bit Mreg218 (Mreg218Out, dataIn, clr, clk, Mreg218Ins);
		reg32bit Mreg219 (Mreg219Out, dataIn, clr, clk, Mreg219Ins);
		reg32bit Mreg220 (Mreg220Out, dataIn, clr, clk, Mreg220Ins);
		reg32bit Mreg221 (Mreg221Out, dataIn, clr, clk, Mreg221Ins);
		reg32bit Mreg222 (Mreg222Out, dataIn, clr, clk, Mreg222Ins);
		reg32bit Mreg223 (Mreg223Out, dataIn, clr, clk, Mreg223Ins);
		reg32bit Mreg224 (Mreg224Out, dataIn, clr, clk, Mreg224Ins);
		reg32bit Mreg225 (Mreg225Out, dataIn, clr, clk, Mreg225Ins);
		reg32bit Mreg226 (Mreg226Out, dataIn, clr, clk, Mreg226Ins);
		reg32bit Mreg227 (Mreg227Out, dataIn, clr, clk, Mreg227Ins);
		reg32bit Mreg228 (Mreg228Out, dataIn, clr, clk, Mreg228Ins);
		reg32bit Mreg229 (Mreg229Out, dataIn, clr, clk, Mreg229Ins);
		reg32bit Mreg230 (Mreg230Out, dataIn, clr, clk, Mreg230Ins);
		reg32bit Mreg231 (Mreg231Out, dataIn, clr, clk, Mreg231Ins);
		reg32bit Mreg232 (Mreg232Out, dataIn, clr, clk, Mreg232Ins);
		reg32bit Mreg233 (Mreg233Out, dataIn, clr, clk, Mreg233Ins);
		reg32bit Mreg234 (Mreg234Out, dataIn, clr, clk, Mreg234Ins);
		reg32bit Mreg235 (Mreg235Out, dataIn, clr, clk, Mreg235Ins);
		reg32bit Mreg236 (Mreg236Out, dataIn, clr, clk, Mreg236Ins);
		reg32bit Mreg237 (Mreg237Out, dataIn, clr, clk, Mreg237Ins);
		reg32bit Mreg238 (Mreg238Out, dataIn, clr, clk, Mreg238Ins);
		reg32bit Mreg239 (Mreg239Out, dataIn, clr, clk, Mreg239Ins);
		reg32bit Mreg240 (Mreg240Out, dataIn, clr, clk, Mreg240Ins);
		reg32bit Mreg241 (Mreg241Out, dataIn, clr, clk, Mreg241Ins);
		reg32bit Mreg242 (Mreg242Out, dataIn, clr, clk, Mreg242Ins);
		reg32bit Mreg243 (Mreg243Out, dataIn, clr, clk, Mreg243Ins);
		reg32bit Mreg244 (Mreg244Out, dataIn, clr, clk, Mreg244Ins);
		reg32bit Mreg245 (Mreg245Out, dataIn, clr, clk, Mreg245Ins);
		reg32bit Mreg246 (Mreg246Out, dataIn, clr, clk, Mreg246Ins);
		reg32bit Mreg247 (Mreg247Out, dataIn, clr, clk, Mreg247Ins);
		reg32bit Mreg248 (Mreg248Out, dataIn, clr, clk, Mreg248Ins);
		reg32bit Mreg249 (Mreg249Out, dataIn, clr, clk, Mreg249Ins);
		reg32bit Mreg250 (Mreg250Out, dataIn, clr, clk, Mreg250Ins);
		reg32bit Mreg251 (Mreg251Out, dataIn, clr, clk, Mreg251Ins);
		reg32bit Mreg252 (Mreg252Out, dataIn, clr, clk, Mreg252Ins);
		reg32bit Mreg253 (Mreg253Out, dataIn, clr, clk, Mreg253Ins);
		reg32bit Mreg254 (Mreg254Out, dataIn, clr, clk, Mreg254Ins);
		reg32bit Mreg255 (Mreg255Out, dataIn, clr, clk, Mreg255Ins);
		reg32bit Mreg256 (Mreg256Out, dataIn, clr, clk, Mreg256Ins);
		reg32bit Mreg257 (Mreg257Out, dataIn, clr, clk, Mreg257Ins);
		reg32bit Mreg258 (Mreg258Out, dataIn, clr, clk, Mreg258Ins);
		reg32bit Mreg259 (Mreg259Out, dataIn, clr, clk, Mreg259Ins);
		reg32bit Mreg260 (Mreg260Out, dataIn, clr, clk, Mreg260Ins);
		reg32bit Mreg261 (Mreg261Out, dataIn, clr, clk, Mreg261Ins);
		reg32bit Mreg262 (Mreg262Out, dataIn, clr, clk, Mreg262Ins);
		reg32bit Mreg263 (Mreg263Out, dataIn, clr, clk, Mreg263Ins);
		reg32bit Mreg264 (Mreg264Out, dataIn, clr, clk, Mreg264Ins);
		reg32bit Mreg265 (Mreg265Out, dataIn, clr, clk, Mreg265Ins);
		reg32bit Mreg266 (Mreg266Out, dataIn, clr, clk, Mreg266Ins);
		reg32bit Mreg267 (Mreg267Out, dataIn, clr, clk, Mreg267Ins);
		reg32bit Mreg268 (Mreg268Out, dataIn, clr, clk, Mreg268Ins);
		reg32bit Mreg269 (Mreg269Out, dataIn, clr, clk, Mreg269Ins);
		reg32bit Mreg270 (Mreg270Out, dataIn, clr, clk, Mreg270Ins);
		reg32bit Mreg271 (Mreg271Out, dataIn, clr, clk, Mreg271Ins);
		reg32bit Mreg272 (Mreg272Out, dataIn, clr, clk, Mreg272Ins);
		reg32bit Mreg273 (Mreg273Out, dataIn, clr, clk, Mreg273Ins);
		reg32bit Mreg274 (Mreg274Out, dataIn, clr, clk, Mreg274Ins);
		reg32bit Mreg275 (Mreg275Out, dataIn, clr, clk, Mreg275Ins);
		reg32bit Mreg276 (Mreg276Out, dataIn, clr, clk, Mreg276Ins);
		reg32bit Mreg277 (Mreg277Out, dataIn, clr, clk, Mreg277Ins);
		reg32bit Mreg278 (Mreg278Out, dataIn, clr, clk, Mreg278Ins);
		reg32bit Mreg279 (Mreg279Out, dataIn, clr, clk, Mreg279Ins);
		reg32bit Mreg280 (Mreg280Out, dataIn, clr, clk, Mreg280Ins);
		reg32bit Mreg281 (Mreg281Out, dataIn, clr, clk, Mreg281Ins);
		reg32bit Mreg282 (Mreg282Out, dataIn, clr, clk, Mreg282Ins);
		reg32bit Mreg283 (Mreg283Out, dataIn, clr, clk, Mreg283Ins);
		reg32bit Mreg284 (Mreg284Out, dataIn, clr, clk, Mreg284Ins);
		reg32bit Mreg285 (Mreg285Out, dataIn, clr, clk, Mreg285Ins);
		reg32bit Mreg286 (Mreg286Out, dataIn, clr, clk, Mreg286Ins);
		reg32bit Mreg287 (Mreg287Out, dataIn, clr, clk, Mreg287Ins);
		reg32bit Mreg288 (Mreg288Out, dataIn, clr, clk, Mreg288Ins);
		reg32bit Mreg289 (Mreg289Out, dataIn, clr, clk, Mreg289Ins);
		reg32bit Mreg290 (Mreg290Out, dataIn, clr, clk, Mreg290Ins);
		reg32bit Mreg291 (Mreg291Out, dataIn, clr, clk, Mreg291Ins);
		reg32bit Mreg292 (Mreg292Out, dataIn, clr, clk, Mreg292Ins);
		reg32bit Mreg293 (Mreg293Out, dataIn, clr, clk, Mreg293Ins);
		reg32bit Mreg294 (Mreg294Out, dataIn, clr, clk, Mreg294Ins);
		reg32bit Mreg295 (Mreg295Out, dataIn, clr, clk, Mreg295Ins);
		reg32bit Mreg296 (Mreg296Out, dataIn, clr, clk, Mreg296Ins);
		reg32bit Mreg297 (Mreg297Out, dataIn, clr, clk, Mreg297Ins);
		reg32bit Mreg298 (Mreg298Out, dataIn, clr, clk, Mreg298Ins);
		reg32bit Mreg299 (Mreg299Out, dataIn, clr, clk, Mreg299Ins);
		//Break for a hundred
		reg32bit Mreg300 (Mreg300Out, dataIn, clr, clk, Mreg300Ins);
		reg32bit Mreg301 (Mreg301Out, dataIn, clr, clk, Mreg301Ins);
		reg32bit Mreg302 (Mreg302Out, dataIn, clr, clk, Mreg302Ins);
		reg32bit Mreg303 (Mreg303Out, dataIn, clr, clk, Mreg303Ins);
		reg32bit Mreg304 (Mreg304Out, dataIn, clr, clk, Mreg304Ins);
		reg32bit Mreg305 (Mreg305Out, dataIn, clr, clk, Mreg305Ins);
		reg32bit Mreg306 (Mreg306Out, dataIn, clr, clk, Mreg306Ins);
		reg32bit Mreg307 (Mreg307Out, dataIn, clr, clk, Mreg307Ins);
		reg32bit Mreg308 (Mreg308Out, dataIn, clr, clk, Mreg308Ins);
		reg32bit Mreg309 (Mreg309Out, dataIn, clr, clk, Mreg309Ins);
		reg32bit Mreg310 (Mreg310Out, dataIn, clr, clk, Mreg310Ins);
		reg32bit Mreg311 (Mreg311Out, dataIn, clr, clk, Mreg311Ins);
		reg32bit Mreg312 (Mreg312Out, dataIn, clr, clk, Mreg312Ins);
		reg32bit Mreg313 (Mreg313Out, dataIn, clr, clk, Mreg313Ins);
		reg32bit Mreg314 (Mreg314Out, dataIn, clr, clk, Mreg314Ins);
		reg32bit Mreg315 (Mreg315Out, dataIn, clr, clk, Mreg315Ins);
		reg32bit Mreg316 (Mreg316Out, dataIn, clr, clk, Mreg316Ins);
		reg32bit Mreg317 (Mreg317Out, dataIn, clr, clk, Mreg317Ins);
		reg32bit Mreg318 (Mreg318Out, dataIn, clr, clk, Mreg318Ins);
		reg32bit Mreg319 (Mreg319Out, dataIn, clr, clk, Mreg319Ins);
		reg32bit Mreg320 (Mreg320Out, dataIn, clr, clk, Mreg320Ins);
		reg32bit Mreg321 (Mreg321Out, dataIn, clr, clk, Mreg321Ins);
		reg32bit Mreg322 (Mreg322Out, dataIn, clr, clk, Mreg322Ins);
		reg32bit Mreg323 (Mreg323Out, dataIn, clr, clk, Mreg323Ins);
		reg32bit Mreg324 (Mreg324Out, dataIn, clr, clk, Mreg324Ins);
		reg32bit Mreg325 (Mreg325Out, dataIn, clr, clk, Mreg325Ins);
		reg32bit Mreg326 (Mreg326Out, dataIn, clr, clk, Mreg326Ins);
		reg32bit Mreg327 (Mreg327Out, dataIn, clr, clk, Mreg327Ins);
		reg32bit Mreg328 (Mreg328Out, dataIn, clr, clk, Mreg328Ins);
		reg32bit Mreg329 (Mreg329Out, dataIn, clr, clk, Mreg329Ins);
		reg32bit Mreg330 (Mreg330Out, dataIn, clr, clk, Mreg330Ins);
		reg32bit Mreg331 (Mreg331Out, dataIn, clr, clk, Mreg331Ins);
		reg32bit Mreg332 (Mreg332Out, dataIn, clr, clk, Mreg332Ins);
		reg32bit Mreg333 (Mreg333Out, dataIn, clr, clk, Mreg333Ins);
		reg32bit Mreg334 (Mreg334Out, dataIn, clr, clk, Mreg334Ins);
		reg32bit Mreg335 (Mreg335Out, dataIn, clr, clk, Mreg335Ins);
		reg32bit Mreg336 (Mreg336Out, dataIn, clr, clk, Mreg336Ins);
		reg32bit Mreg337 (Mreg337Out, dataIn, clr, clk, Mreg337Ins);
		reg32bit Mreg338 (Mreg338Out, dataIn, clr, clk, Mreg338Ins);
		reg32bit Mreg339 (Mreg339Out, dataIn, clr, clk, Mreg339Ins);
		reg32bit Mreg340 (Mreg340Out, dataIn, clr, clk, Mreg340Ins);
		reg32bit Mreg341 (Mreg341Out, dataIn, clr, clk, Mreg341Ins);
		reg32bit Mreg342 (Mreg342Out, dataIn, clr, clk, Mreg342Ins);
		reg32bit Mreg343 (Mreg343Out, dataIn, clr, clk, Mreg343Ins);
		reg32bit Mreg344 (Mreg344Out, dataIn, clr, clk, Mreg344Ins);
		reg32bit Mreg345 (Mreg345Out, dataIn, clr, clk, Mreg345Ins);
		reg32bit Mreg346 (Mreg346Out, dataIn, clr, clk, Mreg346Ins);
		reg32bit Mreg347 (Mreg347Out, dataIn, clr, clk, Mreg347Ins);
		reg32bit Mreg348 (Mreg348Out, dataIn, clr, clk, Mreg348Ins);
		reg32bit Mreg349 (Mreg349Out, dataIn, clr, clk, Mreg349Ins);
		reg32bit Mreg350 (Mreg350Out, dataIn, clr, clk, Mreg350Ins);
		reg32bit Mreg351 (Mreg351Out, dataIn, clr, clk, Mreg351Ins);
		reg32bit Mreg352 (Mreg352Out, dataIn, clr, clk, Mreg352Ins);
		reg32bit Mreg353 (Mreg353Out, dataIn, clr, clk, Mreg353Ins);
		reg32bit Mreg354 (Mreg354Out, dataIn, clr, clk, Mreg354Ins);
		reg32bit Mreg355 (Mreg355Out, dataIn, clr, clk, Mreg355Ins);
		reg32bit Mreg356 (Mreg356Out, dataIn, clr, clk, Mreg356Ins);
		reg32bit Mreg357 (Mreg357Out, dataIn, clr, clk, Mreg357Ins);
		reg32bit Mreg358 (Mreg358Out, dataIn, clr, clk, Mreg358Ins);
		reg32bit Mreg359 (Mreg359Out, dataIn, clr, clk, Mreg359Ins);
		reg32bit Mreg360 (Mreg360Out, dataIn, clr, clk, Mreg360Ins);
		reg32bit Mreg361 (Mreg361Out, dataIn, clr, clk, Mreg361Ins);
		reg32bit Mreg362 (Mreg362Out, dataIn, clr, clk, Mreg362Ins);
		reg32bit Mreg363 (Mreg363Out, dataIn, clr, clk, Mreg363Ins);
		reg32bit Mreg364 (Mreg364Out, dataIn, clr, clk, Mreg364Ins);
		reg32bit Mreg365 (Mreg365Out, dataIn, clr, clk, Mreg365Ins);
		reg32bit Mreg366 (Mreg366Out, dataIn, clr, clk, Mreg366Ins);
		reg32bit Mreg367 (Mreg367Out, dataIn, clr, clk, Mreg367Ins);
		reg32bit Mreg368 (Mreg368Out, dataIn, clr, clk, Mreg368Ins);
		reg32bit Mreg369 (Mreg369Out, dataIn, clr, clk, Mreg369Ins);
		reg32bit Mreg370 (Mreg370Out, dataIn, clr, clk, Mreg370Ins);
		reg32bit Mreg371 (Mreg371Out, dataIn, clr, clk, Mreg371Ins);
		reg32bit Mreg372 (Mreg372Out, dataIn, clr, clk, Mreg372Ins);
		reg32bit Mreg373 (Mreg373Out, dataIn, clr, clk, Mreg373Ins);
		reg32bit Mreg374 (Mreg374Out, dataIn, clr, clk, Mreg374Ins);
		reg32bit Mreg375 (Mreg375Out, dataIn, clr, clk, Mreg375Ins);
		reg32bit Mreg376 (Mreg376Out, dataIn, clr, clk, Mreg376Ins);
		reg32bit Mreg377 (Mreg377Out, dataIn, clr, clk, Mreg377Ins);
		reg32bit Mreg378 (Mreg378Out, dataIn, clr, clk, Mreg378Ins);
		reg32bit Mreg379 (Mreg379Out, dataIn, clr, clk, Mreg379Ins);
		reg32bit Mreg380 (Mreg380Out, dataIn, clr, clk, Mreg380Ins);
		reg32bit Mreg381 (Mreg381Out, dataIn, clr, clk, Mreg381Ins);
		reg32bit Mreg382 (Mreg382Out, dataIn, clr, clk, Mreg382Ins);
		reg32bit Mreg383 (Mreg383Out, dataIn, clr, clk, Mreg383Ins);
		reg32bit Mreg384 (Mreg384Out, dataIn, clr, clk, Mreg384Ins);
		reg32bit Mreg385 (Mreg385Out, dataIn, clr, clk, Mreg385Ins);
		reg32bit Mreg386 (Mreg386Out, dataIn, clr, clk, Mreg386Ins);
		reg32bit Mreg387 (Mreg387Out, dataIn, clr, clk, Mreg387Ins);
		reg32bit Mreg388 (Mreg388Out, dataIn, clr, clk, Mreg388Ins);
		reg32bit Mreg389 (Mreg389Out, dataIn, clr, clk, Mreg389Ins);
		reg32bit Mreg390 (Mreg390Out, dataIn, clr, clk, Mreg390Ins);
		reg32bit Mreg391 (Mreg391Out, dataIn, clr, clk, Mreg391Ins);
		reg32bit Mreg392 (Mreg392Out, dataIn, clr, clk, Mreg392Ins);
		reg32bit Mreg393 (Mreg393Out, dataIn, clr, clk, Mreg393Ins);
		reg32bit Mreg394 (Mreg394Out, dataIn, clr, clk, Mreg394Ins);
		reg32bit Mreg395 (Mreg395Out, dataIn, clr, clk, Mreg395Ins);
		reg32bit Mreg396 (Mreg396Out, dataIn, clr, clk, Mreg396Ins);
		reg32bit Mreg397 (Mreg397Out, dataIn, clr, clk, Mreg397Ins);
		reg32bit Mreg398 (Mreg398Out, dataIn, clr, clk, Mreg398Ins);
		reg32bit Mreg399 (Mreg399Out, dataIn, clr, clk, Mreg399Ins);
		//Break for a hundred
		reg32bit Mreg400 (Mreg400Out, dataIn, clr, clk, Mreg400Ins);
		reg32bit Mreg401 (Mreg401Out, dataIn, clr, clk, Mreg401Ins);
		reg32bit Mreg402 (Mreg402Out, dataIn, clr, clk, Mreg402Ins);
		reg32bit Mreg403 (Mreg403Out, dataIn, clr, clk, Mreg403Ins);
		reg32bit Mreg404 (Mreg404Out, dataIn, clr, clk, Mreg404Ins);
		reg32bit Mreg405 (Mreg405Out, dataIn, clr, clk, Mreg405Ins);
		reg32bit Mreg406 (Mreg406Out, dataIn, clr, clk, Mreg406Ins);
		reg32bit Mreg407 (Mreg407Out, dataIn, clr, clk, Mreg407Ins);
		reg32bit Mreg408 (Mreg408Out, dataIn, clr, clk, Mreg408Ins);
		reg32bit Mreg409 (Mreg409Out, dataIn, clr, clk, Mreg409Ins);
		reg32bit Mreg410 (Mreg410Out, dataIn, clr, clk, Mreg410Ins);
		reg32bit Mreg411 (Mreg411Out, dataIn, clr, clk, Mreg411Ins);
		reg32bit Mreg412 (Mreg412Out, dataIn, clr, clk, Mreg412Ins);
		reg32bit Mreg413 (Mreg413Out, dataIn, clr, clk, Mreg413Ins);
		reg32bit Mreg414 (Mreg414Out, dataIn, clr, clk, Mreg414Ins);
		reg32bit Mreg415 (Mreg415Out, dataIn, clr, clk, Mreg415Ins);
		reg32bit Mreg416 (Mreg416Out, dataIn, clr, clk, Mreg416Ins);
		reg32bit Mreg417 (Mreg417Out, dataIn, clr, clk, Mreg417Ins);
		reg32bit Mreg418 (Mreg418Out, dataIn, clr, clk, Mreg418Ins);
		reg32bit Mreg419 (Mreg419Out, dataIn, clr, clk, Mreg419Ins);
		reg32bit Mreg420 (Mreg420Out, dataIn, clr, clk, Mreg420Ins);
		reg32bit Mreg421 (Mreg421Out, dataIn, clr, clk, Mreg421Ins);
		reg32bit Mreg422 (Mreg422Out, dataIn, clr, clk, Mreg422Ins);
		reg32bit Mreg423 (Mreg423Out, dataIn, clr, clk, Mreg423Ins);
		reg32bit Mreg424 (Mreg424Out, dataIn, clr, clk, Mreg424Ins);
		reg32bit Mreg425 (Mreg425Out, dataIn, clr, clk, Mreg425Ins);
		reg32bit Mreg426 (Mreg426Out, dataIn, clr, clk, Mreg426Ins);
		reg32bit Mreg427 (Mreg427Out, dataIn, clr, clk, Mreg427Ins);
		reg32bit Mreg428 (Mreg428Out, dataIn, clr, clk, Mreg428Ins);
		reg32bit Mreg429 (Mreg429Out, dataIn, clr, clk, Mreg429Ins);
		reg32bit Mreg430 (Mreg430Out, dataIn, clr, clk, Mreg430Ins);
		reg32bit Mreg431 (Mreg431Out, dataIn, clr, clk, Mreg431Ins);
		reg32bit Mreg432 (Mreg432Out, dataIn, clr, clk, Mreg432Ins);
		reg32bit Mreg433 (Mreg433Out, dataIn, clr, clk, Mreg433Ins);
		reg32bit Mreg434 (Mreg434Out, dataIn, clr, clk, Mreg434Ins);
		reg32bit Mreg435 (Mreg435Out, dataIn, clr, clk, Mreg435Ins);
		reg32bit Mreg436 (Mreg436Out, dataIn, clr, clk, Mreg436Ins);
		reg32bit Mreg437 (Mreg437Out, dataIn, clr, clk, Mreg437Ins);
		reg32bit Mreg438 (Mreg438Out, dataIn, clr, clk, Mreg438Ins);
		reg32bit Mreg439 (Mreg439Out, dataIn, clr, clk, Mreg439Ins);
		reg32bit Mreg440 (Mreg440Out, dataIn, clr, clk, Mreg440Ins);
		reg32bit Mreg441 (Mreg441Out, dataIn, clr, clk, Mreg441Ins);
		reg32bit Mreg442 (Mreg442Out, dataIn, clr, clk, Mreg442Ins);
		reg32bit Mreg443 (Mreg443Out, dataIn, clr, clk, Mreg443Ins);
		reg32bit Mreg444 (Mreg444Out, dataIn, clr, clk, Mreg444Ins);
		reg32bit Mreg445 (Mreg445Out, dataIn, clr, clk, Mreg445Ins);
		reg32bit Mreg446 (Mreg446Out, dataIn, clr, clk, Mreg446Ins);
		reg32bit Mreg447 (Mreg447Out, dataIn, clr, clk, Mreg447Ins);
		reg32bit Mreg448 (Mreg448Out, dataIn, clr, clk, Mreg448Ins);
		reg32bit Mreg449 (Mreg449Out, dataIn, clr, clk, Mreg449Ins);
		reg32bit Mreg450 (Mreg450Out, dataIn, clr, clk, Mreg450Ins);
		reg32bit Mreg451 (Mreg451Out, dataIn, clr, clk, Mreg451Ins);
		reg32bit Mreg452 (Mreg452Out, dataIn, clr, clk, Mreg452Ins);
		reg32bit Mreg453 (Mreg453Out, dataIn, clr, clk, Mreg453Ins);
		reg32bit Mreg454 (Mreg454Out, dataIn, clr, clk, Mreg454Ins);
		reg32bit Mreg455 (Mreg455Out, dataIn, clr, clk, Mreg455Ins);
		reg32bit Mreg456 (Mreg456Out, dataIn, clr, clk, Mreg456Ins);
		reg32bit Mreg457 (Mreg457Out, dataIn, clr, clk, Mreg457Ins);
		reg32bit Mreg458 (Mreg458Out, dataIn, clr, clk, Mreg458Ins);
		reg32bit Mreg459 (Mreg459Out, dataIn, clr, clk, Mreg459Ins);
		reg32bit Mreg460 (Mreg460Out, dataIn, clr, clk, Mreg460Ins);
		reg32bit Mreg461 (Mreg461Out, dataIn, clr, clk, Mreg461Ins);
		reg32bit Mreg462 (Mreg462Out, dataIn, clr, clk, Mreg462Ins);
		reg32bit Mreg463 (Mreg463Out, dataIn, clr, clk, Mreg463Ins);
		reg32bit Mreg464 (Mreg464Out, dataIn, clr, clk, Mreg464Ins);
		reg32bit Mreg465 (Mreg465Out, dataIn, clr, clk, Mreg465Ins);
		reg32bit Mreg466 (Mreg466Out, dataIn, clr, clk, Mreg466Ins);
		reg32bit Mreg467 (Mreg467Out, dataIn, clr, clk, Mreg467Ins);
		reg32bit Mreg468 (Mreg468Out, dataIn, clr, clk, Mreg468Ins);
		reg32bit Mreg469 (Mreg469Out, dataIn, clr, clk, Mreg469Ins);
		reg32bit Mreg470 (Mreg470Out, dataIn, clr, clk, Mreg470Ins);
		reg32bit Mreg471 (Mreg471Out, dataIn, clr, clk, Mreg471Ins);
		reg32bit Mreg472 (Mreg472Out, dataIn, clr, clk, Mreg472Ins);
		reg32bit Mreg473 (Mreg473Out, dataIn, clr, clk, Mreg473Ins);
		reg32bit Mreg474 (Mreg474Out, dataIn, clr, clk, Mreg474Ins);
		reg32bit Mreg475 (Mreg475Out, dataIn, clr, clk, Mreg475Ins);
		reg32bit Mreg476 (Mreg476Out, dataIn, clr, clk, Mreg476Ins);
		reg32bit Mreg477 (Mreg477Out, dataIn, clr, clk, Mreg477Ins);
		reg32bit Mreg478 (Mreg478Out, dataIn, clr, clk, Mreg478Ins);
		reg32bit Mreg479 (Mreg479Out, dataIn, clr, clk, Mreg479Ins);
		reg32bit Mreg480 (Mreg480Out, dataIn, clr, clk, Mreg480Ins);
		reg32bit Mreg481 (Mreg481Out, dataIn, clr, clk, Mreg481Ins);
		reg32bit Mreg482 (Mreg482Out, dataIn, clr, clk, Mreg482Ins);
		reg32bit Mreg483 (Mreg483Out, dataIn, clr, clk, Mreg483Ins);
		reg32bit Mreg484 (Mreg484Out, dataIn, clr, clk, Mreg484Ins);
		reg32bit Mreg485 (Mreg485Out, dataIn, clr, clk, Mreg485Ins);
		reg32bit Mreg486 (Mreg486Out, dataIn, clr, clk, Mreg486Ins);
		reg32bit Mreg487 (Mreg487Out, dataIn, clr, clk, Mreg487Ins);
		reg32bit Mreg488 (Mreg488Out, dataIn, clr, clk, Mreg488Ins);
		reg32bit Mreg489 (Mreg489Out, dataIn, clr, clk, Mreg489Ins);
		reg32bit Mreg490 (Mreg490Out, dataIn, clr, clk, Mreg490Ins);
		reg32bit Mreg491 (Mreg491Out, dataIn, clr, clk, Mreg491Ins);
		reg32bit Mreg492 (Mreg492Out, dataIn, clr, clk, Mreg492Ins);
		reg32bit Mreg493 (Mreg493Out, dataIn, clr, clk, Mreg493Ins);
		reg32bit Mreg494 (Mreg494Out, dataIn, clr, clk, Mreg494Ins);
		reg32bit Mreg495 (Mreg495Out, dataIn, clr, clk, Mreg495Ins);
		reg32bit Mreg496 (Mreg496Out, dataIn, clr, clk, Mreg496Ins);
		reg32bit Mreg497 (Mreg497Out, dataIn, clr, clk, Mreg497Ins);
		reg32bit Mreg498 (Mreg498Out, dataIn, clr, clk, Mreg498Ins);
		reg32bit Mreg499 (Mreg499Out, dataIn, clr, clk, Mreg499Ins);
		//Break for a hundred
		reg32bit Mreg500 (Mreg500Out, dataIn, clr, clk, Mreg500Ins);
		reg32bit Mreg501 (Mreg501Out, dataIn, clr, clk, Mreg501Ins);
		reg32bit Mreg502 (Mreg502Out, dataIn, clr, clk, Mreg502Ins);
		reg32bit Mreg503 (Mreg503Out, dataIn, clr, clk, Mreg503Ins);
		reg32bit Mreg504 (Mreg504Out, dataIn, clr, clk, Mreg504Ins);
		reg32bit Mreg505 (Mreg505Out, dataIn, clr, clk, Mreg505Ins);
		reg32bit Mreg506 (Mreg506Out, dataIn, clr, clk, Mreg506Ins);
		reg32bit Mreg507 (Mreg507Out, dataIn, clr, clk, Mreg507Ins);
		reg32bit Mreg508 (Mreg508Out, dataIn, clr, clk, Mreg508Ins);
		reg32bit Mreg509 (Mreg509Out, dataIn, clr, clk, Mreg509Ins);
		reg32bit Mreg510 (Mreg510Out, dataIn, clr, clk, Mreg510Ins);
		reg32bit Mreg511 (Mreg511Out, dataIn, clr, clk, Mreg511Ins);
	endgenerate
	
	//--------------------------------------------------------------------------------------------------------------------------------
	//Finish creation of the registers
	
	//Start the memory write enable decoder
	//--------------------------------------------------------------------------------------------------------------------------------
	always @ (*) begin
		case (Addr)
		9'b000000000 : Mreg0Ins   <= write;
		9'b000000001 : Mreg1Ins   <= write;
		9'b000000010 : Mreg2Ins   <= write;
		9'b000000011 : Mreg3Ins   <= write;
		9'b000000100 : Mreg4Ins   <= write;
		9'b000000101 : Mreg5Ins   <= write;
		9'b000000110 : Mreg6Ins   <= write;
		9'b000000111 : Mreg7Ins   <= write;
		9'b000001000 : Mreg8Ins   <= write;
		9'b000001001 : Mreg9Ins   <= write;
		9'b000001010 : Mreg10Ins  <= write;
		9'b000001011 : Mreg11Ins  <= write;
		9'b000001100 : Mreg12Ins  <= write;
		9'b000001101 : Mreg13Ins  <= write;
		9'b000001110 : Mreg14Ins  <= write;
		9'b000001111 : Mreg15Ins  <= write;
		9'b000010000 : Mreg16Ins  <= write;
		9'b000010001 : Mreg17Ins  <= write;
		9'b000010010 : Mreg18Ins  <= write;
		9'b000010011 : Mreg19Ins  <= write;
		9'b000010100 : Mreg20Ins  <= write;
		9'b000010101 : Mreg21Ins  <= write;
		9'b000010110 : Mreg22Ins  <= write;
		9'b000010111 : Mreg23Ins  <= write;
		9'b000011000 : Mreg24Ins  <= write;
		9'b000011001 : Mreg25Ins  <= write;
		9'b000011010 : Mreg26Ins  <= write;
		9'b000011011 : Mreg27Ins  <= write;
		9'b000011100 : Mreg28Ins  <= write;
		9'b000011101 : Mreg29Ins  <= write;
		9'b000011110 : Mreg30Ins  <= write;
		9'b000011111 : Mreg31Ins  <= write;
		9'b000100000 : Mreg32Ins  <= write;
		9'b000100001 : Mreg33Ins  <= write;
		9'b000100010 : Mreg34Ins  <= write;
		9'b000100011 : Mreg35Ins  <= write;
		9'b000100100 : Mreg36Ins  <= write;
		9'b000100101 : Mreg37Ins  <= write;
		9'b000100110 : Mreg38Ins  <= write;
		9'b000100111 : Mreg39Ins  <= write;
		9'b000101000 : Mreg40Ins  <= write;
		9'b000101001 : Mreg41Ins  <= write;
		9'b000101010 : Mreg42Ins  <= write;
		9'b000101011 : Mreg43Ins  <= write;
		9'b000101100 : Mreg44Ins  <= write;
		9'b000101101 : Mreg45Ins  <= write;
		9'b000101110 : Mreg46Ins  <= write;
		9'b000101111 : Mreg47Ins  <= write;
		9'b000110000 : Mreg48Ins  <= write;
		9'b000110001 : Mreg49Ins  <= write;
		9'b000110010 : Mreg50Ins  <= write;
		9'b000110011 : Mreg51Ins  <= write;
		9'b000110100 : Mreg52Ins  <= write;
		9'b000110101 : Mreg53Ins  <= write;
		9'b000110110 : Mreg54Ins  <= write;
		9'b000110111 : Mreg55Ins  <= write;
		9'b000111000 : Mreg56Ins  <= write;
		9'b000111001 : Mreg57Ins  <= write;
		9'b000111010 : Mreg58Ins  <= write;
		9'b000111011 : Mreg59Ins  <= write;
		9'b000111100 : Mreg60Ins  <= write;
		9'b000111101 : Mreg61Ins  <= write;
		9'b000111110 : Mreg62Ins  <= write;
		9'b000111111 : Mreg63Ins  <= write;
		9'b001000000 : Mreg64Ins  <= write;
		9'b001000001 : Mreg65Ins  <= write;
		9'b001000010 : Mreg66Ins  <= write;
		9'b001000011 : Mreg67Ins  <= write;
		9'b001000100 : Mreg68Ins  <= write;
		9'b001000101 : Mreg69Ins  <= write;
		9'b001000110 : Mreg70Ins  <= write;
		9'b001000111 : Mreg71Ins  <= write;
		9'b001001000 : Mreg72Ins  <= write;
		9'b001001001 : Mreg73Ins  <= write;
		9'b001001010 : Mreg74Ins  <= write;
		9'b001001011 : Mreg75Ins  <= write;
		9'b001001100 : Mreg76Ins  <= write;
		9'b001001101 : Mreg77Ins  <= write;
		9'b001001110 : Mreg78Ins  <= write;
		9'b001001111 : Mreg79Ins  <= write;
		9'b001010000 : Mreg80Ins  <= write;
		9'b001010001 : Mreg81Ins  <= write;
		9'b001010010 : Mreg82Ins  <= write;
		9'b001010011 : Mreg83Ins  <= write;
		9'b001010100 : Mreg84Ins  <= write;
		9'b001010101 : Mreg85Ins  <= write;
		9'b001010110 : Mreg86Ins  <= write;
		9'b001010111 : Mreg87Ins  <= write;
		9'b001011000 : Mreg88Ins  <= write;
		9'b001011001 : Mreg89Ins  <= write;
		9'b001011010 : Mreg90Ins  <= write;
		9'b001011011 : Mreg91Ins  <= write;
		9'b001011100 : Mreg92Ins  <= write;
		9'b001011101 : Mreg93Ins  <= write;
		9'b001011110 : Mreg94Ins  <= write;
		9'b001011111 : Mreg95Ins  <= write;
		9'b001100000 : Mreg96Ins  <= write;
		9'b001100001 : Mreg97Ins  <= write;
		9'b001100010 : Mreg98Ins  <= write;
		9'b001100011 : Mreg99Ins  <= write;
		9'b001100100 : Mreg100Ins <= write;
		9'b001100101 : Mreg101Ins <= write;
		9'b001100110 : Mreg102Ins <= write;
		9'b001100111 : Mreg103Ins <= write;
		9'b001101000 : Mreg104Ins <= write;
		9'b001101001 : Mreg105Ins <= write;
		9'b001101010 : Mreg106Ins <= write;
		9'b001101011 : Mreg107Ins <= write;
		9'b001101100 : Mreg108Ins <= write;
		9'b001101101 : Mreg109Ins <= write;
		9'b001101110 : Mreg110Ins <= write;
		9'b001101111 : Mreg111Ins <= write;
		9'b001110000 : Mreg112Ins <= write;
		9'b001110001 : Mreg113Ins <= write;
		9'b001110010 : Mreg114Ins <= write;
		9'b001110011 : Mreg115Ins <= write;
		9'b001110100 : Mreg116Ins <= write;
		9'b001110101 : Mreg117Ins <= write;
		9'b001110110 : Mreg118Ins <= write;
		9'b001110111 : Mreg119Ins <= write;
		9'b001111000 : Mreg120Ins <= write;
		9'b001111001 : Mreg121Ins <= write;
		9'b001111010 : Mreg122Ins <= write;
		9'b001111011 : Mreg123Ins <= write;
		9'b001111100 : Mreg124Ins <= write;
		9'b001111101 : Mreg125Ins <= write;
		9'b001111110 : Mreg126Ins <= write;
		9'b001111111 : Mreg127Ins <= write;
		9'b010000000 : Mreg128Ins <= write;
		9'b010000001 : Mreg129Ins <= write;
		9'b010000010 : Mreg130Ins <= write;
		9'b010000011 : Mreg131Ins <= write;
		9'b010000100 : Mreg132Ins <= write;
		9'b010000101 : Mreg133Ins <= write;
		9'b010000110 : Mreg134Ins <= write;
		9'b010000111 : Mreg135Ins <= write;
		9'b010001000 : Mreg136Ins <= write;
		9'b010001001 : Mreg137Ins <= write;
		9'b010001010 : Mreg138Ins <= write;
		9'b010001011 : Mreg139Ins <= write;
		9'b010001100 : Mreg140Ins <= write;
		9'b010001101 : Mreg141Ins <= write;
		9'b010001110 : Mreg142Ins <= write;
		9'b010001111 : Mreg143Ins <= write;
		9'b010010000 : Mreg144Ins <= write;
		9'b010010001 : Mreg145Ins <= write;
		9'b010010010 : Mreg146Ins <= write;
		9'b010010011 : Mreg147Ins <= write;
		9'b010010100 : Mreg148Ins <= write;
		9'b010010101 : Mreg149Ins <= write;
		9'b010010110 : Mreg150Ins <= write;
		9'b010010111 : Mreg151Ins <= write;
		9'b010011000 : Mreg152Ins <= write;
		9'b010011001 : Mreg153Ins <= write;
		9'b010011010 : Mreg154Ins <= write;
		9'b010011011 : Mreg155Ins <= write;
		9'b010011100 : Mreg156Ins <= write;
		9'b010011101 : Mreg157Ins <= write;
		9'b010011110 : Mreg158Ins <= write;
		9'b010011111 : Mreg159Ins <= write;
		9'b010100000 : Mreg160Ins <= write;
		9'b010100001 : Mreg161Ins <= write;
		9'b010100010 : Mreg162Ins <= write;
		9'b010100011 : Mreg163Ins <= write;
		9'b010100100 : Mreg164Ins <= write;
		9'b010100101 : Mreg165Ins <= write;
		9'b010100110 : Mreg166Ins <= write;
		9'b010100111 : Mreg167Ins <= write;
		9'b010101000 : Mreg168Ins <= write;
		9'b010101001 : Mreg169Ins <= write;
		9'b010101010 : Mreg170Ins <= write;
		9'b010101011 : Mreg171Ins <= write;
		9'b010101100 : Mreg172Ins <= write;
		9'b010101101 : Mreg173Ins <= write;
		9'b010101110 : Mreg174Ins <= write;
		9'b010101111 : Mreg175Ins <= write;
		9'b010110000 : Mreg176Ins <= write;
		9'b010110001 : Mreg177Ins <= write;
		9'b010110010 : Mreg178Ins <= write;
		9'b010110011 : Mreg179Ins <= write;
		9'b010110100 : Mreg180Ins <= write;
		9'b010110101 : Mreg181Ins <= write;
		9'b010110110 : Mreg182Ins <= write;
		9'b010110111 : Mreg183Ins <= write;
		9'b010111000 : Mreg184Ins <= write;
		9'b010111001 : Mreg185Ins <= write;
		9'b010111010 : Mreg186Ins <= write;
		9'b010111011 : Mreg187Ins <= write;
		9'b010111100 : Mreg188Ins <= write;
		9'b010111101 : Mreg189Ins <= write;
		9'b010111110 : Mreg190Ins <= write;
		9'b010111111 : Mreg191Ins <= write;
		9'b011000000 : Mreg192Ins <= write;
		9'b011000001 : Mreg193Ins <= write;
		9'b011000010 : Mreg194Ins <= write;
		9'b011000011 : Mreg195Ins <= write;
		9'b011000100 : Mreg196Ins <= write;
		9'b011000101 : Mreg197Ins <= write;
		9'b011000110 : Mreg198Ins <= write;
		9'b011000111 : Mreg199Ins <= write;
		9'b011001000 : Mreg200Ins <= write;
		9'b011001001 : Mreg201Ins <= write;
		9'b011001010 : Mreg202Ins <= write;
		9'b011001011 : Mreg203Ins <= write;
		9'b011001100 : Mreg204Ins <= write;
		9'b011001101 : Mreg205Ins <= write;
		9'b011001110 : Mreg206Ins <= write;
		9'b011001111 : Mreg207Ins <= write;
		9'b011010000 : Mreg208Ins <= write;
		9'b011010001 : Mreg209Ins <= write;
		9'b011010010 : Mreg210Ins <= write;
		9'b011010011 : Mreg211Ins <= write;
		9'b011010100 : Mreg212Ins <= write;
		9'b011010101 : Mreg213Ins <= write;
		9'b011010110 : Mreg214Ins <= write;
		9'b011010111 : Mreg215Ins <= write;
		9'b011011000 : Mreg216Ins <= write;
		9'b011011001 : Mreg217Ins <= write;
		9'b011011010 : Mreg218Ins <= write;
		9'b011011011 : Mreg219Ins <= write;
		9'b011011100 : Mreg220Ins <= write;
		9'b011011101 : Mreg221Ins <= write;
		9'b011011110 : Mreg222Ins <= write;
		9'b011011111 : Mreg223Ins <= write;
		9'b011100000 : Mreg224Ins <= write;
		9'b011100001 : Mreg225Ins <= write;
		9'b011100010 : Mreg226Ins <= write;
		9'b011100011 : Mreg227Ins <= write;
		9'b011100100 : Mreg228Ins <= write;
		9'b011100101 : Mreg229Ins <= write;
		9'b011100110 : Mreg230Ins <= write;
		9'b011100111 : Mreg231Ins <= write;
		9'b011101000 : Mreg232Ins <= write;
		9'b011101001 : Mreg233Ins <= write;
		9'b011101010 : Mreg234Ins <= write;
		9'b011101011 : Mreg235Ins <= write;
		9'b011101100 : Mreg236Ins <= write;
		9'b011101101 : Mreg237Ins <= write;
		9'b011101110 : Mreg238Ins <= write;
		9'b011101111 : Mreg239Ins <= write;
		9'b011110000 : Mreg240Ins <= write;
		9'b011110001 : Mreg241Ins <= write;
		9'b011110010 : Mreg242Ins <= write;
		9'b011110011 : Mreg243Ins <= write;
		9'b011110100 : Mreg244Ins <= write;
		9'b011110101 : Mreg245Ins <= write;
		9'b011110110 : Mreg246Ins <= write;
		9'b011110111 : Mreg247Ins <= write;
		9'b011111000 : Mreg248Ins <= write;
		9'b011111001 : Mreg249Ins <= write;
		9'b011111010 : Mreg250Ins <= write;
		9'b011111011 : Mreg251Ins <= write;
		9'b011111100 : Mreg252Ins <= write;
		9'b011111101 : Mreg253Ins <= write;
		9'b011111110 : Mreg254Ins <= write;
		9'b011111111 : Mreg255Ins <= write;
		9'b100000000 : Mreg256Ins <= write;
		9'b100000001 : Mreg257Ins <= write;
		9'b100000010 : Mreg258Ins <= write;
		9'b100000011 : Mreg259Ins <= write;
		9'b100000100 : Mreg260Ins <= write;
		9'b100000101 : Mreg261Ins <= write;
		9'b100000110 : Mreg262Ins <= write;
		9'b100000111 : Mreg263Ins <= write;
		9'b100001000 : Mreg264Ins <= write;
		9'b100001001 : Mreg265Ins <= write;
		9'b100001010 : Mreg266Ins <= write;
		9'b100001011 : Mreg267Ins <= write;
		9'b100001100 : Mreg268Ins <= write;
		9'b100001101 : Mreg269Ins <= write;
		9'b100001110 : Mreg270Ins <= write;
		9'b100001111 : Mreg271Ins <= write;
		9'b100010000 : Mreg272Ins <= write;
		9'b100010001 : Mreg273Ins <= write;
		9'b100010010 : Mreg274Ins <= write;
		9'b100010011 : Mreg275Ins <= write;
		9'b100010100 : Mreg276Ins <= write;
		9'b100010101 : Mreg277Ins <= write;
		9'b100010110 : Mreg278Ins <= write;
		9'b100010111 : Mreg279Ins <= write;
		9'b100011000 : Mreg280Ins <= write;
		9'b100011001 : Mreg281Ins <= write;
		9'b100011010 : Mreg282Ins <= write;
		9'b100011011 : Mreg283Ins <= write;
		9'b100011100 : Mreg284Ins <= write;
		9'b100011101 : Mreg285Ins <= write;
		9'b100011110 : Mreg286Ins <= write;
		9'b100011111 : Mreg287Ins <= write;
		9'b100100000 : Mreg288Ins <= write;
		9'b100100001 : Mreg289Ins <= write;
		9'b100100010 : Mreg290Ins <= write;
		9'b100100011 : Mreg291Ins <= write;
		9'b100100100 : Mreg292Ins <= write;
		9'b100100101 : Mreg293Ins <= write;
		9'b100100110 : Mreg294Ins <= write;
		9'b100100111 : Mreg295Ins <= write;
		9'b100101000 : Mreg296Ins <= write;
		9'b100101001 : Mreg297Ins <= write;
		9'b100101010 : Mreg298Ins <= write;
		9'b100101011 : Mreg299Ins <= write;
		9'b100101100 : Mreg300Ins <= write;
		9'b100101101 : Mreg301Ins <= write;
		9'b100101110 : Mreg302Ins <= write;
		9'b100101111 : Mreg303Ins <= write;
		9'b100110000 : Mreg304Ins <= write;
		9'b100110001 : Mreg305Ins <= write;
		9'b100110010 : Mreg306Ins <= write;
		9'b100110011 : Mreg307Ins <= write;
		9'b100110100 : Mreg308Ins <= write;
		9'b100110101 : Mreg309Ins <= write;
		9'b100110110 : Mreg310Ins <= write;
		9'b100110111 : Mreg311Ins <= write;
		9'b100111000 : Mreg312Ins <= write;
		9'b100111001 : Mreg313Ins <= write;
		9'b100111010 : Mreg314Ins <= write;
		9'b100111011 : Mreg315Ins <= write;
		9'b100111100 : Mreg316Ins <= write;
		9'b100111101 : Mreg317Ins <= write;
		9'b100111110 : Mreg318Ins <= write;
		9'b100111111 : Mreg319Ins <= write;
		9'b101000000 : Mreg320Ins <= write;
		9'b101000001 : Mreg321Ins <= write;
		9'b101000010 : Mreg322Ins <= write;
		9'b101000011 : Mreg323Ins <= write;
		9'b101000100 : Mreg324Ins <= write;
		9'b101000101 : Mreg325Ins <= write;
		9'b101000110 : Mreg326Ins <= write;
		9'b101000111 : Mreg327Ins <= write;
		9'b101001000 : Mreg328Ins <= write;
		9'b101001001 : Mreg329Ins <= write;
		9'b101001010 : Mreg330Ins <= write;
		9'b101001011 : Mreg331Ins <= write;
		9'b101001100 : Mreg332Ins <= write;
		9'b101001101 : Mreg333Ins <= write;
		9'b101001110 : Mreg334Ins <= write;
		9'b101001111 : Mreg335Ins <= write;
		9'b101010000 : Mreg336Ins <= write;
		9'b101010001 : Mreg337Ins <= write;
		9'b101010010 : Mreg338Ins <= write;
		9'b101010011 : Mreg339Ins <= write;
		9'b101010100 : Mreg340Ins <= write;
		9'b101010101 : Mreg341Ins <= write;
		9'b101010110 : Mreg342Ins <= write;
		9'b101010111 : Mreg343Ins <= write;
		9'b101011000 : Mreg344Ins <= write;
		9'b101011001 : Mreg345Ins <= write;
		9'b101011010 : Mreg346Ins <= write;
		9'b101011011 : Mreg347Ins <= write;
		9'b101011100 : Mreg348Ins <= write;
		9'b101011101 : Mreg349Ins <= write;
		9'b101011110 : Mreg350Ins <= write;
		9'b101011111 : Mreg351Ins <= write;
		9'b101100000 : Mreg352Ins <= write;
		9'b101100001 : Mreg353Ins <= write;
		9'b101100010 : Mreg354Ins <= write;
		9'b101100011 : Mreg355Ins <= write;
		9'b101100100 : Mreg356Ins <= write;
		9'b101100101 : Mreg357Ins <= write;
		9'b101100110 : Mreg358Ins <= write;
		9'b101100111 : Mreg359Ins <= write;
		9'b101101000 : Mreg360Ins <= write;
		9'b101101001 : Mreg361Ins <= write;
		9'b101101010 : Mreg362Ins <= write;
		9'b101101011 : Mreg363Ins <= write;
		9'b101101100 : Mreg364Ins <= write;
		9'b101101101 : Mreg365Ins <= write;
		9'b101101110 : Mreg366Ins <= write;
		9'b101101111 : Mreg367Ins <= write;
		9'b101110000 : Mreg368Ins <= write;
		9'b101110001 : Mreg369Ins <= write;
		9'b101110010 : Mreg370Ins <= write;
		9'b101110011 : Mreg371Ins <= write;
		9'b101110100 : Mreg372Ins <= write;
		9'b101110101 : Mreg373Ins <= write;
		9'b101110110 : Mreg374Ins <= write;
		9'b101110111 : Mreg375Ins <= write;
		9'b101111000 : Mreg376Ins <= write;
		9'b101111001 : Mreg377Ins <= write;
		9'b101111010 : Mreg378Ins <= write;
		9'b101111011 : Mreg379Ins <= write;
		9'b101111100 : Mreg380Ins <= write;
		9'b101111101 : Mreg381Ins <= write;
		9'b101111110 : Mreg382Ins <= write;
		9'b101111111 : Mreg383Ins <= write;
		9'b110000000 : Mreg384Ins <= write;
		9'b110000001 : Mreg385Ins <= write;
		9'b110000010 : Mreg386Ins <= write;
		9'b110000011 : Mreg387Ins <= write;
		9'b110000100 : Mreg388Ins <= write;
		9'b110000101 : Mreg389Ins <= write;
		9'b110000110 : Mreg390Ins <= write;
		9'b110000111 : Mreg391Ins <= write;
		9'b110001000 : Mreg392Ins <= write;
		9'b110001001 : Mreg393Ins <= write;
		9'b110001010 : Mreg394Ins <= write;
		9'b110001011 : Mreg395Ins <= write;
		9'b110001100 : Mreg396Ins <= write;
		9'b110001101 : Mreg397Ins <= write;
		9'b110001110 : Mreg398Ins <= write;
		9'b110001111 : Mreg399Ins <= write;
		9'b110010000 : Mreg400Ins <= write;
		9'b110010001 : Mreg401Ins <= write;
		9'b110010010 : Mreg402Ins <= write;
		9'b110010011 : Mreg403Ins <= write;
		9'b110010100 : Mreg404Ins <= write;
		9'b110010101 : Mreg405Ins <= write;
		9'b110010110 : Mreg406Ins <= write;
		9'b110010111 : Mreg407Ins <= write;
		9'b110011000 : Mreg408Ins <= write;
		9'b110011001 : Mreg409Ins <= write;
		9'b110011010 : Mreg410Ins <= write;
		9'b110011011 : Mreg411Ins <= write;
		9'b110011100 : Mreg412Ins <= write;
		9'b110011101 : Mreg413Ins <= write;
		9'b110011110 : Mreg414Ins <= write;
		9'b110011111 : Mreg415Ins <= write;
		9'b110100000 : Mreg416Ins <= write;
		9'b110100001 : Mreg417Ins <= write;
		9'b110100010 : Mreg418Ins <= write;
		9'b110100011 : Mreg419Ins <= write;
		9'b110100100 : Mreg420Ins <= write;
		9'b110100101 : Mreg421Ins <= write;
		9'b110100110 : Mreg422Ins <= write;
		9'b110100111 : Mreg423Ins <= write;
		9'b110101000 : Mreg424Ins <= write;
		9'b110101001 : Mreg425Ins <= write;
		9'b110101010 : Mreg426Ins <= write;
		9'b110101011 : Mreg427Ins <= write;
		9'b110101100 : Mreg428Ins <= write;
		9'b110101101 : Mreg429Ins <= write;
		9'b110101110 : Mreg430Ins <= write;
		9'b110101111 : Mreg431Ins <= write;
		9'b110110000 : Mreg432Ins <= write;
		9'b110110001 : Mreg433Ins <= write;
		9'b110110010 : Mreg434Ins <= write;
		9'b110110011 : Mreg435Ins <= write;
		9'b110110100 : Mreg436Ins <= write;
		9'b110110101 : Mreg437Ins <= write;
		9'b110110110 : Mreg438Ins <= write;
		9'b110110111 : Mreg439Ins <= write;
		9'b110111000 : Mreg440Ins <= write;
		9'b110111001 : Mreg441Ins <= write;
		9'b110111010 : Mreg442Ins <= write;
		9'b110111011 : Mreg443Ins <= write;
		9'b110111100 : Mreg444Ins <= write;
		9'b110111101 : Mreg445Ins <= write;
		9'b110111110 : Mreg446Ins <= write;
		9'b110111111 : Mreg447Ins <= write;
		9'b111000000 : Mreg448Ins <= write;
		9'b111000001 : Mreg449Ins <= write;
		9'b111000010 : Mreg450Ins <= write;
		9'b111000011 : Mreg451Ins <= write;
		9'b111000100 : Mreg452Ins <= write;
		9'b111000101 : Mreg453Ins <= write;
		9'b111000110 : Mreg454Ins <= write;
		9'b111000111 : Mreg455Ins <= write;
		9'b111001000 : Mreg456Ins <= write;
		9'b111001001 : Mreg457Ins <= write;
		9'b111001010 : Mreg458Ins <= write;
		9'b111001011 : Mreg459Ins <= write;
		9'b111001100 : Mreg460Ins <= write;
		9'b111001101 : Mreg461Ins <= write;
		9'b111001110 : Mreg462Ins <= write;
		9'b111001111 : Mreg463Ins <= write;
		9'b111010000 : Mreg464Ins <= write;
		9'b111010001 : Mreg465Ins <= write;
		9'b111010010 : Mreg466Ins <= write;
		9'b111010011 : Mreg467Ins <= write;
		9'b111010100 : Mreg468Ins <= write;
		9'b111010101 : Mreg469Ins <= write;
		9'b111010110 : Mreg470Ins <= write;
		9'b111010111 : Mreg471Ins <= write;
		9'b111011000 : Mreg472Ins <= write;
		9'b111011001 : Mreg473Ins <= write;
		9'b111011010 : Mreg474Ins <= write;
		9'b111011011 : Mreg475Ins <= write;
		9'b111011100 : Mreg476Ins <= write;
		9'b111011101 : Mreg477Ins <= write;
		9'b111011110 : Mreg478Ins <= write;
		9'b111011111 : Mreg479Ins <= write;
		9'b111100000 : Mreg480Ins <= write;
		9'b111100001 : Mreg481Ins <= write;
		9'b111100010 : Mreg482Ins <= write;
		9'b111100011 : Mreg483Ins <= write;
		9'b111100100 : Mreg484Ins <= write;
		9'b111100101 : Mreg485Ins <= write;
		9'b111100110 : Mreg486Ins <= write;
		9'b111100111 : Mreg487Ins <= write;
		9'b111101000 : Mreg488Ins <= write;
		9'b111101001 : Mreg489Ins <= write;
		9'b111101010 : Mreg490Ins <= write;
		9'b111101011 : Mreg491Ins <= write;
		9'b111101100 : Mreg492Ins <= write;
		9'b111101101 : Mreg493Ins <= write;
		9'b111101110 : Mreg494Ins <= write;
		9'b111101111 : Mreg495Ins <= write;
		9'b111110000 : Mreg496Ins <= write;
		9'b111110001 : Mreg497Ins <= write;
		9'b111110010 : Mreg498Ins <= write;
		9'b111110011 : Mreg499Ins <= write;
		9'b111110100 : Mreg500Ins <= write;
		9'b111110101 : Mreg501Ins <= write;
		9'b111110110 : Mreg502Ins <= write;
		9'b111110111 : Mreg503Ins <= write;
		9'b111111000 : Mreg504Ins <= write;
		9'b111111001 : Mreg505Ins <= write;
		9'b111111010 : Mreg506Ins <= write;
		9'b111111011 : Mreg507Ins <= write;
		9'b111111100 : Mreg508Ins <= write;
		9'b111111101 : Mreg509Ins <= write;
		9'b111111110 : Mreg510Ins <= write;
		9'b111111111 : Mreg511Ins <= write; 
	endcase	
end
	//--------------------------------------------------------------------------------------------------------------------------------
	//Finish the memory write enable decoder
	
	//Start the memory output multiplexer
	//--------------------------------------------------------------------------------------------------------------------------------
	always @ (*) begin
		case (Addr)
		9'b000000000 : dataOutTemp <= Mreg0Out  ; 
		9'b000000001 : dataOutTemp <= Mreg1Out  ; 
		9'b000000010 : dataOutTemp <= Mreg2Out  ; 
		9'b000000011 : dataOutTemp <= Mreg3Out  ; 
		9'b000000100 : dataOutTemp <= Mreg4Out  ; 
		9'b000000101 : dataOutTemp <= Mreg5Out  ; 
		9'b000000110 : dataOutTemp <= Mreg6Out  ; 
		9'b000000111 : dataOutTemp <= Mreg7Out  ; 
		9'b000001000 : dataOutTemp <= Mreg8Out  ; 
		9'b000001001 : dataOutTemp <= Mreg9Out  ; 
		9'b000001010 : dataOutTemp <= Mreg10Out ; 
		9'b000001011 : dataOutTemp <= Mreg11Out ; 
		9'b000001100 : dataOutTemp <= Mreg12Out ; 
		9'b000001101 : dataOutTemp <= Mreg13Out ; 
		9'b000001110 : dataOutTemp <= Mreg14Out ; 
		9'b000001111 : dataOutTemp <= Mreg15Out ; 
		9'b000010000 : dataOutTemp <= Mreg16Out ; 
		9'b000010001 : dataOutTemp <= Mreg17Out ; 
		9'b000010010 : dataOutTemp <= Mreg18Out ; 
		9'b000010011 : dataOutTemp <= Mreg19Out ; 
		9'b000010100 : dataOutTemp <= Mreg20Out ; 
		9'b000010101 : dataOutTemp <= Mreg21Out ; 
		9'b000010110 : dataOutTemp <= Mreg22Out ; 
		9'b000010111 : dataOutTemp <= Mreg23Out ; 
		9'b000011000 : dataOutTemp <= Mreg24Out ; 
		9'b000011001 : dataOutTemp <= Mreg25Out ; 
		9'b000011010 : dataOutTemp <= Mreg26Out ; 
		9'b000011011 : dataOutTemp <= Mreg27Out ; 
		9'b000011100 : dataOutTemp <= Mreg28Out ; 
		9'b000011101 : dataOutTemp <= Mreg29Out ; 
		9'b000011110 : dataOutTemp <= Mreg30Out ; 
		9'b000011111 : dataOutTemp <= Mreg31Out ; 
		9'b000100000 : dataOutTemp <= Mreg32Out ; 
		9'b000100001 : dataOutTemp <= Mreg33Out ; 
		9'b000100010 : dataOutTemp <= Mreg34Out ; 
		9'b000100011 : dataOutTemp <= Mreg35Out ; 
		9'b000100100 : dataOutTemp <= Mreg36Out ; 
		9'b000100101 : dataOutTemp <= Mreg37Out ; 
		9'b000100110 : dataOutTemp <= Mreg38Out ; 
		9'b000100111 : dataOutTemp <= Mreg39Out ; 
		9'b000101000 : dataOutTemp <= Mreg40Out ; 
		9'b000101001 : dataOutTemp <= Mreg41Out ; 
		9'b000101010 : dataOutTemp <= Mreg42Out ; 
		9'b000101011 : dataOutTemp <= Mreg43Out ; 
		9'b000101100 : dataOutTemp <= Mreg44Out ; 
		9'b000101101 : dataOutTemp <= Mreg45Out ; 
		9'b000101110 : dataOutTemp <= Mreg46Out ; 
		9'b000101111 : dataOutTemp <= Mreg47Out ; 
		9'b000110000 : dataOutTemp <= Mreg48Out ; 
		9'b000110001 : dataOutTemp <= Mreg49Out ; 
		9'b000110010 : dataOutTemp <= Mreg50Out ; 
		9'b000110011 : dataOutTemp <= Mreg51Out ; 
		9'b000110100 : dataOutTemp <= Mreg52Out ; 
		9'b000110101 : dataOutTemp <= Mreg53Out ; 
		9'b000110110 : dataOutTemp <= Mreg54Out ; 
		9'b000110111 : dataOutTemp <= Mreg55Out ; 
		9'b000111000 : dataOutTemp <= Mreg56Out ; 
		9'b000111001 : dataOutTemp <= Mreg57Out ; 
		9'b000111010 : dataOutTemp <= Mreg58Out ; 
		9'b000111011 : dataOutTemp <= Mreg59Out ; 
		9'b000111100 : dataOutTemp <= Mreg60Out ; 
		9'b000111101 : dataOutTemp <= Mreg61Out ; 
		9'b000111110 : dataOutTemp <= Mreg62Out ; 
		9'b000111111 : dataOutTemp <= Mreg63Out ; 
		9'b001000000 : dataOutTemp <= Mreg64Out ; 
		9'b001000001 : dataOutTemp <= Mreg65Out ; 
		9'b001000010 : dataOutTemp <= Mreg66Out ; 
		9'b001000011 : dataOutTemp <= Mreg67Out ; 
		9'b001000100 : dataOutTemp <= Mreg68Out ; 
		9'b001000101 : dataOutTemp <= Mreg69Out ; 
		9'b001000110 : dataOutTemp <= Mreg70Out ; 
		9'b001000111 : dataOutTemp <= Mreg71Out ; 
		9'b001001000 : dataOutTemp <= Mreg72Out ; 
		9'b001001001 : dataOutTemp <= Mreg73Out ; 
		9'b001001010 : dataOutTemp <= Mreg74Out ; 
		9'b001001011 : dataOutTemp <= Mreg75Out ; 
		9'b001001100 : dataOutTemp <= Mreg76Out ; 
		9'b001001101 : dataOutTemp <= Mreg77Out ; 
		9'b001001110 : dataOutTemp <= Mreg78Out ; 
		9'b001001111 : dataOutTemp <= Mreg79Out ; 
		9'b001010000 : dataOutTemp <= Mreg80Out ; 
		9'b001010001 : dataOutTemp <= Mreg81Out ; 
		9'b001010010 : dataOutTemp <= Mreg82Out ; 
		9'b001010011 : dataOutTemp <= Mreg83Out ; 
		9'b001010100 : dataOutTemp <= Mreg84Out ; 
		9'b001010101 : dataOutTemp <= Mreg85Out ; 
		9'b001010110 : dataOutTemp <= Mreg86Out ; 
		9'b001010111 : dataOutTemp <= Mreg87Out ; 
		9'b001011000 : dataOutTemp <= Mreg88Out ; 
		9'b001011001 : dataOutTemp <= Mreg89Out ; 
		9'b001011010 : dataOutTemp <= Mreg90Out ; 
		9'b001011011 : dataOutTemp <= Mreg91Out ; 
		9'b001011100 : dataOutTemp <= Mreg92Out ; 
		9'b001011101 : dataOutTemp <= Mreg93Out ; 
		9'b001011110 : dataOutTemp <= Mreg94Out ; 
		9'b001011111 : dataOutTemp <= Mreg95Out ; 
		9'b001100000 : dataOutTemp <= Mreg96Out ; 
		9'b001100001 : dataOutTemp <= Mreg97Out ; 
		9'b001100010 : dataOutTemp <= Mreg98Out ; 
		9'b001100011 : dataOutTemp <= Mreg99Out ; 
		9'b001100100 : dataOutTemp <= Mreg100Out; 
		9'b001100101 : dataOutTemp <= Mreg101Out; 
		9'b001100110 : dataOutTemp <= Mreg102Out; 
		9'b001100111 : dataOutTemp <= Mreg103Out; 
		9'b001101000 : dataOutTemp <= Mreg104Out; 
		9'b001101001 : dataOutTemp <= Mreg105Out; 
		9'b001101010 : dataOutTemp <= Mreg106Out; 
		9'b001101011 : dataOutTemp <= Mreg107Out; 
		9'b001101100 : dataOutTemp <= Mreg108Out; 
		9'b001101101 : dataOutTemp <= Mreg109Out; 
		9'b001101110 : dataOutTemp <= Mreg110Out; 
		9'b001101111 : dataOutTemp <= Mreg111Out; 
		9'b001110000 : dataOutTemp <= Mreg112Out; 
		9'b001110001 : dataOutTemp <= Mreg113Out; 
		9'b001110010 : dataOutTemp <= Mreg114Out; 
		9'b001110011 : dataOutTemp <= Mreg115Out; 
		9'b001110100 : dataOutTemp <= Mreg116Out; 
		9'b001110101 : dataOutTemp <= Mreg117Out; 
		9'b001110110 : dataOutTemp <= Mreg118Out; 
		9'b001110111 : dataOutTemp <= Mreg119Out; 
		9'b001111000 : dataOutTemp <= Mreg120Out; 
		9'b001111001 : dataOutTemp <= Mreg121Out; 
		9'b001111010 : dataOutTemp <= Mreg122Out; 
		9'b001111011 : dataOutTemp <= Mreg123Out; 
		9'b001111100 : dataOutTemp <= Mreg124Out; 
		9'b001111101 : dataOutTemp <= Mreg125Out; 
		9'b001111110 : dataOutTemp <= Mreg126Out; 
		9'b001111111 : dataOutTemp <= Mreg127Out; 
		9'b010000000 : dataOutTemp <= Mreg128Out; 
		9'b010000001 : dataOutTemp <= Mreg129Out; 
		9'b010000010 : dataOutTemp <= Mreg130Out; 
		9'b010000011 : dataOutTemp <= Mreg131Out; 
		9'b010000100 : dataOutTemp <= Mreg132Out; 
		9'b010000101 : dataOutTemp <= Mreg133Out; 
		9'b010000110 : dataOutTemp <= Mreg134Out; 
		9'b010000111 : dataOutTemp <= Mreg135Out; 
		9'b010001000 : dataOutTemp <= Mreg136Out; 
		9'b010001001 : dataOutTemp <= Mreg137Out; 
		9'b010001010 : dataOutTemp <= Mreg138Out; 
		9'b010001011 : dataOutTemp <= Mreg139Out; 
		9'b010001100 : dataOutTemp <= Mreg140Out; 
		9'b010001101 : dataOutTemp <= Mreg141Out; 
		9'b010001110 : dataOutTemp <= Mreg142Out; 
		9'b010001111 : dataOutTemp <= Mreg143Out; 
		9'b010010000 : dataOutTemp <= Mreg144Out; 
		9'b010010001 : dataOutTemp <= Mreg145Out; 
		9'b010010010 : dataOutTemp <= Mreg146Out; 
		9'b010010011 : dataOutTemp <= Mreg147Out; 
		9'b010010100 : dataOutTemp <= Mreg148Out; 
		9'b010010101 : dataOutTemp <= Mreg149Out; 
		9'b010010110 : dataOutTemp <= Mreg150Out; 
		9'b010010111 : dataOutTemp <= Mreg151Out; 
		9'b010011000 : dataOutTemp <= Mreg152Out; 
		9'b010011001 : dataOutTemp <= Mreg153Out; 
		9'b010011010 : dataOutTemp <= Mreg154Out; 
		9'b010011011 : dataOutTemp <= Mreg155Out; 
		9'b010011100 : dataOutTemp <= Mreg156Out; 
		9'b010011101 : dataOutTemp <= Mreg157Out; 
		9'b010011110 : dataOutTemp <= Mreg158Out; 
		9'b010011111 : dataOutTemp <= Mreg159Out; 
		9'b010100000 : dataOutTemp <= Mreg160Out; 
		9'b010100001 : dataOutTemp <= Mreg161Out; 
		9'b010100010 : dataOutTemp <= Mreg162Out; 
		9'b010100011 : dataOutTemp <= Mreg163Out; 
		9'b010100100 : dataOutTemp <= Mreg164Out; 
		9'b010100101 : dataOutTemp <= Mreg165Out; 
		9'b010100110 : dataOutTemp <= Mreg166Out; 
		9'b010100111 : dataOutTemp <= Mreg167Out; 
		9'b010101000 : dataOutTemp <= Mreg168Out; 
		9'b010101001 : dataOutTemp <= Mreg169Out; 
		9'b010101010 : dataOutTemp <= Mreg170Out; 
		9'b010101011 : dataOutTemp <= Mreg171Out; 
		9'b010101100 : dataOutTemp <= Mreg172Out; 
		9'b010101101 : dataOutTemp <= Mreg173Out; 
		9'b010101110 : dataOutTemp <= Mreg174Out; 
		9'b010101111 : dataOutTemp <= Mreg175Out; 
		9'b010110000 : dataOutTemp <= Mreg176Out; 
		9'b010110001 : dataOutTemp <= Mreg177Out; 
		9'b010110010 : dataOutTemp <= Mreg178Out; 
		9'b010110011 : dataOutTemp <= Mreg179Out; 
		9'b010110100 : dataOutTemp <= Mreg180Out; 
		9'b010110101 : dataOutTemp <= Mreg181Out; 
		9'b010110110 : dataOutTemp <= Mreg182Out; 
		9'b010110111 : dataOutTemp <= Mreg183Out; 
		9'b010111000 : dataOutTemp <= Mreg184Out; 
		9'b010111001 : dataOutTemp <= Mreg185Out; 
		9'b010111010 : dataOutTemp <= Mreg186Out; 
		9'b010111011 : dataOutTemp <= Mreg187Out; 
		9'b010111100 : dataOutTemp <= Mreg188Out; 
		9'b010111101 : dataOutTemp <= Mreg189Out; 
		9'b010111110 : dataOutTemp <= Mreg190Out; 
		9'b010111111 : dataOutTemp <= Mreg191Out; 
		9'b011000000 : dataOutTemp <= Mreg192Out; 
		9'b011000001 : dataOutTemp <= Mreg193Out; 
		9'b011000010 : dataOutTemp <= Mreg194Out; 
		9'b011000011 : dataOutTemp <= Mreg195Out; 
		9'b011000100 : dataOutTemp <= Mreg196Out; 
		9'b011000101 : dataOutTemp <= Mreg197Out; 
		9'b011000110 : dataOutTemp <= Mreg198Out; 
		9'b011000111 : dataOutTemp <= Mreg199Out; 
		9'b011001000 : dataOutTemp <= Mreg200Out; 
		9'b011001001 : dataOutTemp <= Mreg201Out; 
		9'b011001010 : dataOutTemp <= Mreg202Out; 
		9'b011001011 : dataOutTemp <= Mreg203Out; 
		9'b011001100 : dataOutTemp <= Mreg204Out; 
		9'b011001101 : dataOutTemp <= Mreg205Out; 
		9'b011001110 : dataOutTemp <= Mreg206Out; 
		9'b011001111 : dataOutTemp <= Mreg207Out; 
		9'b011010000 : dataOutTemp <= Mreg208Out; 
		9'b011010001 : dataOutTemp <= Mreg209Out; 
		9'b011010010 : dataOutTemp <= Mreg210Out; 
		9'b011010011 : dataOutTemp <= Mreg211Out; 
		9'b011010100 : dataOutTemp <= Mreg212Out; 
		9'b011010101 : dataOutTemp <= Mreg213Out; 
		9'b011010110 : dataOutTemp <= Mreg214Out; 
		9'b011010111 : dataOutTemp <= Mreg215Out; 
		9'b011011000 : dataOutTemp <= Mreg216Out; 
		9'b011011001 : dataOutTemp <= Mreg217Out; 
		9'b011011010 : dataOutTemp <= Mreg218Out; 
		9'b011011011 : dataOutTemp <= Mreg219Out; 
		9'b011011100 : dataOutTemp <= Mreg220Out; 
		9'b011011101 : dataOutTemp <= Mreg221Out; 
		9'b011011110 : dataOutTemp <= Mreg222Out; 
		9'b011011111 : dataOutTemp <= Mreg223Out; 
		9'b011100000 : dataOutTemp <= Mreg224Out; 
		9'b011100001 : dataOutTemp <= Mreg225Out; 
		9'b011100010 : dataOutTemp <= Mreg226Out; 
		9'b011100011 : dataOutTemp <= Mreg227Out; 
		9'b011100100 : dataOutTemp <= Mreg228Out; 
		9'b011100101 : dataOutTemp <= Mreg229Out; 
		9'b011100110 : dataOutTemp <= Mreg230Out; 
		9'b011100111 : dataOutTemp <= Mreg231Out; 
		9'b011101000 : dataOutTemp <= Mreg232Out; 
		9'b011101001 : dataOutTemp <= Mreg233Out; 
		9'b011101010 : dataOutTemp <= Mreg234Out; 
		9'b011101011 : dataOutTemp <= Mreg235Out; 
		9'b011101100 : dataOutTemp <= Mreg236Out; 
		9'b011101101 : dataOutTemp <= Mreg237Out; 
		9'b011101110 : dataOutTemp <= Mreg238Out; 
		9'b011101111 : dataOutTemp <= Mreg239Out; 
		9'b011110000 : dataOutTemp <= Mreg240Out; 
		9'b011110001 : dataOutTemp <= Mreg241Out; 
		9'b011110010 : dataOutTemp <= Mreg242Out; 
		9'b011110011 : dataOutTemp <= Mreg243Out; 
		9'b011110100 : dataOutTemp <= Mreg244Out; 
		9'b011110101 : dataOutTemp <= Mreg245Out; 
		9'b011110110 : dataOutTemp <= Mreg246Out; 
		9'b011110111 : dataOutTemp <= Mreg247Out; 
		9'b011111000 : dataOutTemp <= Mreg248Out; 
		9'b011111001 : dataOutTemp <= Mreg249Out; 
		9'b011111010 : dataOutTemp <= Mreg250Out; 
		9'b011111011 : dataOutTemp <= Mreg251Out; 
		9'b011111100 : dataOutTemp <= Mreg252Out; 
		9'b011111101 : dataOutTemp <= Mreg253Out; 
		9'b011111110 : dataOutTemp <= Mreg254Out; 
		9'b011111111 : dataOutTemp <= Mreg255Out; 
		9'b100000000 : dataOutTemp <= Mreg256Out; 
		9'b100000001 : dataOutTemp <= Mreg257Out; 
		9'b100000010 : dataOutTemp <= Mreg258Out; 
		9'b100000011 : dataOutTemp <= Mreg259Out; 
		9'b100000100 : dataOutTemp <= Mreg260Out; 
		9'b100000101 : dataOutTemp <= Mreg261Out; 
		9'b100000110 : dataOutTemp <= Mreg262Out; 
		9'b100000111 : dataOutTemp <= Mreg263Out; 
		9'b100001000 : dataOutTemp <= Mreg264Out; 
		9'b100001001 : dataOutTemp <= Mreg265Out; 
		9'b100001010 : dataOutTemp <= Mreg266Out; 
		9'b100001011 : dataOutTemp <= Mreg267Out; 
		9'b100001100 : dataOutTemp <= Mreg268Out; 
		9'b100001101 : dataOutTemp <= Mreg269Out; 
		9'b100001110 : dataOutTemp <= Mreg270Out; 
		9'b100001111 : dataOutTemp <= Mreg271Out; 
		9'b100010000 : dataOutTemp <= Mreg272Out; 
		9'b100010001 : dataOutTemp <= Mreg273Out; 
		9'b100010010 : dataOutTemp <= Mreg274Out; 
		9'b100010011 : dataOutTemp <= Mreg275Out; 
		9'b100010100 : dataOutTemp <= Mreg276Out; 
		9'b100010101 : dataOutTemp <= Mreg277Out; 
		9'b100010110 : dataOutTemp <= Mreg278Out; 
		9'b100010111 : dataOutTemp <= Mreg279Out; 
		9'b100011000 : dataOutTemp <= Mreg280Out; 
		9'b100011001 : dataOutTemp <= Mreg281Out; 
		9'b100011010 : dataOutTemp <= Mreg282Out; 
		9'b100011011 : dataOutTemp <= Mreg283Out; 
		9'b100011100 : dataOutTemp <= Mreg284Out; 
		9'b100011101 : dataOutTemp <= Mreg285Out; 
		9'b100011110 : dataOutTemp <= Mreg286Out; 
		9'b100011111 : dataOutTemp <= Mreg287Out; 
		9'b100100000 : dataOutTemp <= Mreg288Out; 
		9'b100100001 : dataOutTemp <= Mreg289Out; 
		9'b100100010 : dataOutTemp <= Mreg290Out; 
		9'b100100011 : dataOutTemp <= Mreg291Out; 
		9'b100100100 : dataOutTemp <= Mreg292Out; 
		9'b100100101 : dataOutTemp <= Mreg293Out; 
		9'b100100110 : dataOutTemp <= Mreg294Out; 
		9'b100100111 : dataOutTemp <= Mreg295Out; 
		9'b100101000 : dataOutTemp <= Mreg296Out; 
		9'b100101001 : dataOutTemp <= Mreg297Out; 
		9'b100101010 : dataOutTemp <= Mreg298Out; 
		9'b100101011 : dataOutTemp <= Mreg299Out; 
		9'b100101100 : dataOutTemp <= Mreg300Out; 
		9'b100101101 : dataOutTemp <= Mreg301Out; 
		9'b100101110 : dataOutTemp <= Mreg302Out; 
		9'b100101111 : dataOutTemp <= Mreg303Out; 
		9'b100110000 : dataOutTemp <= Mreg304Out; 
		9'b100110001 : dataOutTemp <= Mreg305Out; 
		9'b100110010 : dataOutTemp <= Mreg306Out; 
		9'b100110011 : dataOutTemp <= Mreg307Out; 
		9'b100110100 : dataOutTemp <= Mreg308Out; 
		9'b100110101 : dataOutTemp <= Mreg309Out; 
		9'b100110110 : dataOutTemp <= Mreg310Out; 
		9'b100110111 : dataOutTemp <= Mreg311Out; 
		9'b100111000 : dataOutTemp <= Mreg312Out; 
		9'b100111001 : dataOutTemp <= Mreg313Out; 
		9'b100111010 : dataOutTemp <= Mreg314Out; 
		9'b100111011 : dataOutTemp <= Mreg315Out; 
		9'b100111100 : dataOutTemp <= Mreg316Out; 
		9'b100111101 : dataOutTemp <= Mreg317Out; 
		9'b100111110 : dataOutTemp <= Mreg318Out; 
		9'b100111111 : dataOutTemp <= Mreg319Out; 
		9'b101000000 : dataOutTemp <= Mreg320Out; 
		9'b101000001 : dataOutTemp <= Mreg321Out; 
		9'b101000010 : dataOutTemp <= Mreg322Out; 
		9'b101000011 : dataOutTemp <= Mreg323Out; 
		9'b101000100 : dataOutTemp <= Mreg324Out; 
		9'b101000101 : dataOutTemp <= Mreg325Out; 
		9'b101000110 : dataOutTemp <= Mreg326Out; 
		9'b101000111 : dataOutTemp <= Mreg327Out; 
		9'b101001000 : dataOutTemp <= Mreg328Out; 
		9'b101001001 : dataOutTemp <= Mreg329Out; 
		9'b101001010 : dataOutTemp <= Mreg330Out; 
		9'b101001011 : dataOutTemp <= Mreg331Out; 
		9'b101001100 : dataOutTemp <= Mreg332Out; 
		9'b101001101 : dataOutTemp <= Mreg333Out; 
		9'b101001110 : dataOutTemp <= Mreg334Out; 
		9'b101001111 : dataOutTemp <= Mreg335Out; 
		9'b101010000 : dataOutTemp <= Mreg336Out; 
		9'b101010001 : dataOutTemp <= Mreg337Out; 
		9'b101010010 : dataOutTemp <= Mreg338Out; 
		9'b101010011 : dataOutTemp <= Mreg339Out; 
		9'b101010100 : dataOutTemp <= Mreg340Out; 
		9'b101010101 : dataOutTemp <= Mreg341Out; 
		9'b101010110 : dataOutTemp <= Mreg342Out; 
		9'b101010111 : dataOutTemp <= Mreg343Out; 
		9'b101011000 : dataOutTemp <= Mreg344Out; 
		9'b101011001 : dataOutTemp <= Mreg345Out; 
		9'b101011010 : dataOutTemp <= Mreg346Out; 
		9'b101011011 : dataOutTemp <= Mreg347Out; 
		9'b101011100 : dataOutTemp <= Mreg348Out; 
		9'b101011101 : dataOutTemp <= Mreg349Out; 
		9'b101011110 : dataOutTemp <= Mreg350Out; 
		9'b101011111 : dataOutTemp <= Mreg351Out; 
		9'b101100000 : dataOutTemp <= Mreg352Out; 
		9'b101100001 : dataOutTemp <= Mreg353Out; 
		9'b101100010 : dataOutTemp <= Mreg354Out; 
		9'b101100011 : dataOutTemp <= Mreg355Out; 
		9'b101100100 : dataOutTemp <= Mreg356Out; 
		9'b101100101 : dataOutTemp <= Mreg357Out; 
		9'b101100110 : dataOutTemp <= Mreg358Out; 
		9'b101100111 : dataOutTemp <= Mreg359Out; 
		9'b101101000 : dataOutTemp <= Mreg360Out; 
		9'b101101001 : dataOutTemp <= Mreg361Out; 
		9'b101101010 : dataOutTemp <= Mreg362Out; 
		9'b101101011 : dataOutTemp <= Mreg363Out; 
		9'b101101100 : dataOutTemp <= Mreg364Out; 
		9'b101101101 : dataOutTemp <= Mreg365Out; 
		9'b101101110 : dataOutTemp <= Mreg366Out; 
		9'b101101111 : dataOutTemp <= Mreg367Out; 
		9'b101110000 : dataOutTemp <= Mreg368Out; 
		9'b101110001 : dataOutTemp <= Mreg369Out; 
		9'b101110010 : dataOutTemp <= Mreg370Out; 
		9'b101110011 : dataOutTemp <= Mreg371Out; 
		9'b101110100 : dataOutTemp <= Mreg372Out; 
		9'b101110101 : dataOutTemp <= Mreg373Out; 
		9'b101110110 : dataOutTemp <= Mreg374Out; 
		9'b101110111 : dataOutTemp <= Mreg375Out; 
		9'b101111000 : dataOutTemp <= Mreg376Out; 
		9'b101111001 : dataOutTemp <= Mreg377Out; 
		9'b101111010 : dataOutTemp <= Mreg378Out; 
		9'b101111011 : dataOutTemp <= Mreg379Out; 
		9'b101111100 : dataOutTemp <= Mreg380Out; 
		9'b101111101 : dataOutTemp <= Mreg381Out; 
		9'b101111110 : dataOutTemp <= Mreg382Out; 
		9'b101111111 : dataOutTemp <= Mreg383Out; 
		9'b110000000 : dataOutTemp <= Mreg384Out; 
		9'b110000001 : dataOutTemp <= Mreg385Out; 
		9'b110000010 : dataOutTemp <= Mreg386Out; 
		9'b110000011 : dataOutTemp <= Mreg387Out; 
		9'b110000100 : dataOutTemp <= Mreg388Out; 
		9'b110000101 : dataOutTemp <= Mreg389Out; 
		9'b110000110 : dataOutTemp <= Mreg390Out; 
		9'b110000111 : dataOutTemp <= Mreg391Out; 
		9'b110001000 : dataOutTemp <= Mreg392Out; 
		9'b110001001 : dataOutTemp <= Mreg393Out; 
		9'b110001010 : dataOutTemp <= Mreg394Out; 
		9'b110001011 : dataOutTemp <= Mreg395Out; 
		9'b110001100 : dataOutTemp <= Mreg396Out; 
		9'b110001101 : dataOutTemp <= Mreg397Out; 
		9'b110001110 : dataOutTemp <= Mreg398Out; 
		9'b110001111 : dataOutTemp <= Mreg399Out; 
		9'b110010000 : dataOutTemp <= Mreg400Out; 
		9'b110010001 : dataOutTemp <= Mreg401Out; 
		9'b110010010 : dataOutTemp <= Mreg402Out; 
		9'b110010011 : dataOutTemp <= Mreg403Out; 
		9'b110010100 : dataOutTemp <= Mreg404Out; 
		9'b110010101 : dataOutTemp <= Mreg405Out; 
		9'b110010110 : dataOutTemp <= Mreg406Out; 
		9'b110010111 : dataOutTemp <= Mreg407Out; 
		9'b110011000 : dataOutTemp <= Mreg408Out; 
		9'b110011001 : dataOutTemp <= Mreg409Out; 
		9'b110011010 : dataOutTemp <= Mreg410Out; 
		9'b110011011 : dataOutTemp <= Mreg411Out; 
		9'b110011100 : dataOutTemp <= Mreg412Out; 
		9'b110011101 : dataOutTemp <= Mreg413Out; 
		9'b110011110 : dataOutTemp <= Mreg414Out; 
		9'b110011111 : dataOutTemp <= Mreg415Out; 
		9'b110100000 : dataOutTemp <= Mreg416Out; 
		9'b110100001 : dataOutTemp <= Mreg417Out; 
		9'b110100010 : dataOutTemp <= Mreg418Out; 
		9'b110100011 : dataOutTemp <= Mreg419Out; 
		9'b110100100 : dataOutTemp <= Mreg420Out; 
		9'b110100101 : dataOutTemp <= Mreg421Out; 
		9'b110100110 : dataOutTemp <= Mreg422Out; 
		9'b110100111 : dataOutTemp <= Mreg423Out; 
		9'b110101000 : dataOutTemp <= Mreg424Out; 
		9'b110101001 : dataOutTemp <= Mreg425Out; 
		9'b110101010 : dataOutTemp <= Mreg426Out; 
		9'b110101011 : dataOutTemp <= Mreg427Out; 
		9'b110101100 : dataOutTemp <= Mreg428Out; 
		9'b110101101 : dataOutTemp <= Mreg429Out; 
		9'b110101110 : dataOutTemp <= Mreg430Out; 
		9'b110101111 : dataOutTemp <= Mreg431Out; 
		9'b110110000 : dataOutTemp <= Mreg432Out; 
		9'b110110001 : dataOutTemp <= Mreg433Out; 
		9'b110110010 : dataOutTemp <= Mreg434Out; 
		9'b110110011 : dataOutTemp <= Mreg435Out; 
		9'b110110100 : dataOutTemp <= Mreg436Out; 
		9'b110110101 : dataOutTemp <= Mreg437Out; 
		9'b110110110 : dataOutTemp <= Mreg438Out; 
		9'b110110111 : dataOutTemp <= Mreg439Out; 
		9'b110111000 : dataOutTemp <= Mreg440Out; 
		9'b110111001 : dataOutTemp <= Mreg441Out; 
		9'b110111010 : dataOutTemp <= Mreg442Out; 
		9'b110111011 : dataOutTemp <= Mreg443Out; 
		9'b110111100 : dataOutTemp <= Mreg444Out; 
		9'b110111101 : dataOutTemp <= Mreg445Out; 
		9'b110111110 : dataOutTemp <= Mreg446Out; 
		9'b110111111 : dataOutTemp <= Mreg447Out; 
		9'b111000000 : dataOutTemp <= Mreg448Out; 
		9'b111000001 : dataOutTemp <= Mreg449Out; 
		9'b111000010 : dataOutTemp <= Mreg450Out; 
		9'b111000011 : dataOutTemp <= Mreg451Out; 
		9'b111000100 : dataOutTemp <= Mreg452Out; 
		9'b111000101 : dataOutTemp <= Mreg453Out; 
		9'b111000110 : dataOutTemp <= Mreg454Out; 
		9'b111000111 : dataOutTemp <= Mreg455Out; 
		9'b111001000 : dataOutTemp <= Mreg456Out; 
		9'b111001001 : dataOutTemp <= Mreg457Out; 
		9'b111001010 : dataOutTemp <= Mreg458Out; 
		9'b111001011 : dataOutTemp <= Mreg459Out; 
		9'b111001100 : dataOutTemp <= Mreg460Out; 
		9'b111001101 : dataOutTemp <= Mreg461Out; 
		9'b111001110 : dataOutTemp <= Mreg462Out; 
		9'b111001111 : dataOutTemp <= Mreg463Out; 
		9'b111010000 : dataOutTemp <= Mreg464Out; 
		9'b111010001 : dataOutTemp <= Mreg465Out; 
		9'b111010010 : dataOutTemp <= Mreg466Out; 
		9'b111010011 : dataOutTemp <= Mreg467Out; 
		9'b111010100 : dataOutTemp <= Mreg468Out; 
		9'b111010101 : dataOutTemp <= Mreg469Out; 
		9'b111010110 : dataOutTemp <= Mreg470Out; 
		9'b111010111 : dataOutTemp <= Mreg471Out; 
		9'b111011000 : dataOutTemp <= Mreg472Out; 
		9'b111011001 : dataOutTemp <= Mreg473Out; 
		9'b111011010 : dataOutTemp <= Mreg474Out; 
		9'b111011011 : dataOutTemp <= Mreg475Out; 
		9'b111011100 : dataOutTemp <= Mreg476Out; 
		9'b111011101 : dataOutTemp <= Mreg477Out; 
		9'b111011110 : dataOutTemp <= Mreg478Out; 
		9'b111011111 : dataOutTemp <= Mreg479Out; 
		9'b111100000 : dataOutTemp <= Mreg480Out; 
		9'b111100001 : dataOutTemp <= Mreg481Out; 
		9'b111100010 : dataOutTemp <= Mreg482Out; 
		9'b111100011 : dataOutTemp <= Mreg483Out; 
		9'b111100100 : dataOutTemp <= Mreg484Out; 
		9'b111100101 : dataOutTemp <= Mreg485Out; 
		9'b111100110 : dataOutTemp <= Mreg486Out; 
		9'b111100111 : dataOutTemp <= Mreg487Out; 
		9'b111101000 : dataOutTemp <= Mreg488Out; 
		9'b111101001 : dataOutTemp <= Mreg489Out; 
		9'b111101010 : dataOutTemp <= Mreg490Out; 
		9'b111101011 : dataOutTemp <= Mreg491Out; 
		9'b111101100 : dataOutTemp <= Mreg492Out; 
		9'b111101101 : dataOutTemp <= Mreg493Out; 
		9'b111101110 : dataOutTemp <= Mreg494Out; 
		9'b111101111 : dataOutTemp <= Mreg495Out; 
		9'b111110000 : dataOutTemp <= Mreg496Out; 
		9'b111110001 : dataOutTemp <= Mreg497Out; 
		9'b111110010 : dataOutTemp <= Mreg498Out; 
		9'b111110011 : dataOutTemp <= Mreg499Out; 
		9'b111110100 : dataOutTemp <= Mreg500Out; 
		9'b111110101 : dataOutTemp <= Mreg501Out; 
		9'b111110110 : dataOutTemp <= Mreg502Out; 
		9'b111110111 : dataOutTemp <= Mreg503Out; 
		9'b111111000 : dataOutTemp <= Mreg504Out; 
		9'b111111001 : dataOutTemp <= Mreg505Out; 
		9'b111111010 : dataOutTemp <= Mreg506Out; 
		9'b111111011 : dataOutTemp <= Mreg507Out; 
		9'b111111100 : dataOutTemp <= Mreg508Out; 
		9'b111111101 : dataOutTemp <= Mreg509Out; 
		9'b111111110 : dataOutTemp <= Mreg510Out; 
		9'b111111111 : dataOutTemp <= Mreg511Out; 
	endcase
end
	//--------------------------------------------------------------------------------------------------------------------------------
	//Finish the memory output multiplexer
	
assign dataOut = dataOutTemp;
endmodule 